��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���麍�Ks�%$����+d7��/��������ߔ,���<�E�]��&��z>��>�X�����`��B�㓪F:��ew���@�C�k�.U6�vά1�xrl9��Sr?$R�t��M��~3pwd��<�i��w_�)4ޟo$#)����4F�1s[�p;��Q�!����7�5G��Ξ@��/6����=;+�Cgt�ܫ����ߥo��yqa�ĝ!�G�F#{5� �E؃��\il����A�E�sƸ��]��i��Y���i���	��'i�6�9U�x� ��n���}FA3Yt��SRJ��UZ��	����\�\�t[�oA��g��m�o�I��뚑	�u�!y7� С��/wn�31h�O�3�8w|?���oh��m�&��}���Af�m*tH��i�U����W��-�JһS����si���Z�v�x�謙���FMW�K$��r��R����-�OMjK>I4H��;�}�������brQ0�݋1,
�TSt�Kh?u	�,`���i7���3����J{UMÂ�sA҆�z?|�~�x��5�D��Ę�w�]����g�}��.�|���O9A�n�L����f�D��m �ds{��3.�Z�?��' �u�]�L(�����g!�Y���FAW��� ��q�;Wy9w�Q�! ��5����h��O�w8̜*��9{a^W
�����@�AM�FEd�,~Ū�Xm0o�B��'q�_%�fQ���l�k��/��\�g6g���`�Hb���s��o�k+z�L��|;�b��*���{��7&OKZr�}�W��I��*ξ������� X��a.sޗ�Zx�8Xp�?!S�*1"$���^�j�B�J�<�.��1"��ˁs}�J�*�1Z�w�����
���T&T����dJ!զ�>Y���q���ݤ��c5��c�}��V>��p�i*Y���,�����夹SA{�Ǡr���:޸��S�>��(��R����}��;rT��ZwsR���Z��|�m�00���4B|�`�i�>����+?N���6�93|����Zl�� �����kZ�%�|;)<��4˪c2��g��.��3������>��!��9����H�Q"^n��i��3F�Y��n�4^9�B+ҶHp��0jr�
_��Pu]s#YX��.��+�-���l�=���o)��	ev�#���'$�����S���{ɴ��Pκވ��<[���P	�����X�J���A���	ev���~�Nw���E�C܈k��͞��5A(Sa�G&0�{L*e|C����%S�f+�S��NRW�|�� ������:��f�"��C���;�e��K����@�mÈ`=�zV��OȒ�:�y	!��I�g�j�^��'#F�#綏0 $�H���������n�������x2N��H  CVg���:4�Z�d��>��K����u�z����
u9h�eVekuqE4A��=f��� ���B����hW5��8�?~��qa�'���Nf
1�pI�/T��vmK/�f\#��E�	h��~Ff��:������f���s�\�3d����y���)��2L5H�m�?f��!]����Ǌ��iR:��$|mRFt���&%߯.���о�`�]�`��г�]T��c���7�zԶ�]X�}de�����Ȭ~pI�O��T{�Tb�"ń�̢{�px�}et�Щn���,o��2�$�}��d74_�R�)����c\����<^��]f_b�Y�E��V� ����G���}�')�"WQ/��!�R�Gr�׹Ea<�1���'R���pɟ����W����TS��0xJ�i�|�9�L`�.ٞ4z��«�Cj�(��Q��G���uE���i�Ϸ��CUR�
�j�+?�k�m1M���S�7�(=!�-�{�h���!/.da��e�9��^�B���-��dR�cS����$\M_�H�����P�<'���U�m�޻z-��iċ���������(f�7Ԛ'��ӣ�E��C�-]��Oz�� ;�A���o���\$�=��g����l�T+�b��[u�i��H22�ʂ����?\�M<���L,L,���>�]=���CБ�6�x���,64����U5%-�$]P�0����aӐ������ѩ=�Нă�Ml�I�7�/ca�y�˞o�<�d02�[�������������|�)���;���#H�=(�q��#��:�4���H��JU��F>c�����8qV�����!'ξ2���o���H<b8�����W�;sZex��k�b�é�jg�%���F>7ūFBv|�^�*�=���U)�o}Xg͎g	o�2�Kt�岳aB�aY�^�ދM�g��x�C��]Y��.u�乵N
��G �is��j$��vG$0V�9�ߡsaA�w�H�_��[���{/�<����xKi�� ��y��ƀfё���+:�l�	�fz�"��5�%q�
��F�RD�ҵ�O,���i����a<�;l��0�$���%
�eՅ�U��U���Y��	Z�W���+�8[�L>';��)V�l�Z1�s��9�~3���m,/$�����@̣6�#X�B	5H�s��}���H%�9�px����ׄ��6���Ew?'yϜ��-kbb�e��3�����9\Y�ChbhS�w�����ՙ�-b|H�h�q�2w�8R��R/>
ʹ�N�S�~�sz����G����0�;�2� �%7N���Y�qx�c�x5&��;��'֧<f�U�8���'��f�D̊����"���r*{/�v��g:�9cpP�}H�%1Gt���[WH*�=����̊���RŘ�u��E���U�,�~O�Q�U���}jC?
���࡯��B ���gi�x�`<�[�FiUV�C��1�o3Lgd Ų2'�������F�13��Å3���b8/{f@���8�`�ܼ�9�R��~Bbo`>w�%\�q�\��X�^@<�o�Y�o���E _Uq���u9x�pE����A#}c�6d1;�Xz�y��-֫{�O�M��a�Cl�K�)�#�R~q��K��ަ������eέ��z�.���w��K�#~#N\�_��d��D5�`�x�U��f� _�Y_s��� ��3��H8��3���@̈́:�(d��8�/G@x:�N^%��� Wx���^�FJ���k���F�)T����H�}��=c�v�^�a�/
�]�c�GsE\8�Nӌ�.(e�'�x^dZ�l�v��8�_���	1tC��Oէ;dp�2���S�?�|+y��w�P���76>`�l���8In�-�����s�@��r �Y$2*��qO��͌����<IN�KT���s�E��kQ�^80��2^S��si�j��"eM+���E�U�KQ��4`s��w���&܈[���3]!0;��֔��%�!Q�9�}Q]�9���#�.��!%'�)@�x��	�K3� 鈫J]��� o���_�8�崀�I����w��Z�,y�4�evFԂ��UoC�zcj��Y3O�sG���Ոo���q�NV!��+
�%�dkݶ������S�K/�`L(�tZ(S��Ğ�f�\y�8�W~�����Y���R�о�q���?9D��z�I6������!QnC-�Da��x[��]�Ə��[a������ɋG�&}*�뿤����L��5��vM:!���{���"U�t�d�yX�\g�PZ��j�X��h���Q@9�˫b�5�xx%y�{���E�I?�Cĭr;���~X\�4�vr���Ÿ��q�Ҭ��E1�;B}g����rf�Ҧ��
����@��E�t_B�L�=j���,�2��`�+ ;@���)N�?ִ�1W���h��Ul%t@)���o�y����
�Ll�E4�,��e�h��;���I��\y(tQ�d��m�R��{�����A��KT�_NV!�Htt��)KP��J��L�'JY�FB���,ay�;|�o׳���F��nk',t(j֩�09��zhk�8�b�Mrw�c+��⨭�e!�	h@c�Ug�v��Kۃ�d��⪡�a�7i� j�[�O����e��w��ה�UX��A��Mo!XP���{Ԑ��Z��k8�Qe��L>����:�a%1���J�z�W��/���+C��c�o[�p��b���z�# �Ūd���b: �����be����n�#[�じ�![ID�R�S�m�gR���JS�4SKR�gz���3zf��[ܭg���=cue�aަ�\ey+�Rw�H�����X�Ӧ���i�p g聾1����J���U-<h�Q7~�%�p'��D/��=�0S���5eY��%5?	uQ�0S���O��_F���}H�MJ#�������c]��;�nm�ҁ��j��!Q���܎�;�R�04��oߝ��QKKo��9�W~�n��n���R�H}Ԃ]��b�[w��z����>tzݼ����RjL�f��j2�ue����N�'�@��0U��n�S�W&e�<�3ڴ�e���ƕz�I �[7����q{E%c=oC5.����2���F����\U>���d3������ǧ���꥖{�Q����r3���+!6XPU��n;��'�1_�ǈ��Gr;A�*4��;�%*�.��ʬ��-0N�C�p��$ݼ@�7��H� �)a����AI���=,6�kŐ>Ub�����eB�� ����)�:tm��B	�K�f��oF����X>]]�	7:�'�JS?�>��LK'�����/�߈:��Zk<J�|����A��J}w�-b�}w�����-��DK�_����1[:N�?�Q�߫�n��jZ=1�:Nf��J��SĹ�<R�]֧��xu�W�O�O���V�~��%��N%C��LO��z�2�tI!�7�{��g���D"r� � �K:lF����X?&��vZԪ��%չ�d^gZ�ͦ�Ԑ��|��J���jK�^�ZbL���`}�4k}��~�ؔ7��(h��c�)����,��6���`������?����:�V��<���N����J徵r� �Yt4,r��ǯ=K����l��&�6pdS4e�U}d�U�s�����Jr:LS��K46� W������K� <�8��ט7;)o���{�W�YŮR �S0�@�NE�'j�2��'m֢����Cc<��E��9��0�_��G�p�3�^��f+%��f|Iz��Y
���>����m�G����vM��_�E_ Ř��m�-�睻o]1�Ϳ2:,�j�T�s�Q��?�j�mP3=�;>��D4�	t��+��P��>�~g�R�C��H���N�ь�4��1�R�����4��?�P"h����i�.fe�P��)���X��0�L���HJB��rKi�{aR~S�Z��
�koo� 7��� @\�ӯ�l��x��7�/i��@��p ���><]C�_��	�l.#�X����;kτ�gx��ux�J�hD�X1��	78��gN3��>x�A^Oۇ�ɌoS�G�60�l���S�>�Y�"�Gu�/m���ܢ�б}|jE϶�Z��g��b� ՟���D������6W�An�-!Pʋ
+�GӋ}U��@@�km������D�n8)��U�Z��m�9����Ϡ�>X�'�uF��s�&��`=O����~K�7ش32�f��x� �Vv��~\T]�s�K������?��a���uL���C���u�@Bl��c�
�4m�)���L��g��^'V K��KWm��ޡ�B�0o=��7�-�HE��t�Iҗ� ����v`��7��5�,�5���z`	��
���k1&�{[!*v?Q9��+:f���?OFl�;'Z?h]
Tx����G����Dq
OD�*H�n��+��v:8,��T2�T&����Su�lL��Xej�j�/Kl6s��?ĻzF��F�a�YO��6dZ�OS��S��W��*U�ؤX�	�O-�_�D�D�m�$b�����x@�Mce�zX�So�=R�Pa�ύ�����Zq���`礼�x����+0vI*Z}��P7n����4+��`,�"���q=�L��ݜH���i�$'Y�ӧ���R�a��3�Uŉ��. Q>������=���K�M�^�ݱړc���"�ꢗ�</v>�ȎPo�iV^�O��?~�;Y*�ͫ7['0�0���|j��v�nV��	N��q�x� ����ԇ���;$�i,L���;^}H� ���7K2���4��!w���_-ݥĥ�*0�
��h�L�(�z��$i0�R<�6�;�o��L	v�:>X�n��op��G��?N�!Z�ZƊ��ٺ���ͥ�۪9��:k���U������i`�Mj��bN	��8�������������,�c?��2�A�_����\WvJ�I���}mƸ�g3f�g�ʢ�_	C����V�'6 �� Yp����r&���Uچi��Bw�L���k�q�o�O	i���+�����|jW\� h,�@P��B�/5��A�|,ԺU��P�_
͹oc�H�Y����LO�^�կ96�'������Ώljƿo��=�o`�p�-}��/��Y���v�k��+�,��/̿������!�DdC��r6jǵ^/0���J)�>�<��m9�O�r>q���#N�Q�E� ;�� f0z�rB�>y��La�~���7{�af��>�5�����u'�'ˑb�U���$��yu	 UR{5����0zj�{�� �k���{H�VW�X,ʢ,-2[{s�C⤧�C�1oȌ�χ�*�����ٵ�\c�
J|"aiQ��v�����EĸWƹ;�F>o]a��Sd<7$�*kt%�=d���pʃ�OU<��r��0[c׬�f��N�'��ժ�A���c�t%Ps�M��	ƙ.��G}�GM^@9��;ך�V��2�x�>*Έ�j�N~/O.��~����i��o��Ֆ"(\��ED2:*�o}1�lZݛ]�.�k��4wE��c��?�����F�o4�xs���=�rE��6�S08�|*����AxѲ�̾�C�ln�#�K�Iy�l�:�p�҇�V��X�����+�����\W�c��A5>(�"R�9x��?�cKEU���u`�%��F����>'�����/+V��P�0��a0�z�$�q��!� d���M��e���z��f��)'p��N�G�4L��7c₹%�3(W��~Bu�̍��i(��(̾PWY��OH͓4��3��B^�ҫѤ�E�fW�*�Xަ���!���WE�ݲ��R�{_�N�A���I?a9�����/B��
����<hAٛ��jӁ0����i�w�ܝ�i+�yއ�U[\k�F줼�j�h�� U���H��#�}��Hpn��*�ⅾ%�s^:��,WD�Ų�x���L�n A�@ :i޻�h���/�@�t]��v��w2;��uT�C�v���4=x��'�"C��0B�3-\�%{�����e�ls���Q_�� h,^�7���������iS`ֱ���4��0����������p(�
H�c�}���c�`qW\h
9}r�����Tk�(��݇Y�54��������m�;/X'��J#O��J[B�P�w^���t�Ѭ*1h2�ÃYyE��9�����t�2��������D:^�c�u��5a���\i ��'�>;�KG�Ԕ���c(�n[���m��F��s	>E{�:3�8ڋ�����c�H|z����H��r?q�Y'����^��\t������}���(O3��}|v2w��������F��W�4���cF1�v�H�R�s~�*��շ+��5��i��v52����07ݛh�	ٲ�WK�!���_m!�<�J���ײ(������Hp��l�+j������8{�@aV��\�8��d�&ZQƶ�W���m=E�/O��� ���=��v3'I����Mx*��D#�H�tD��s�E�<����Gf����)y�W�����������w��PZ;�f�&��4����M�d=<����g��f�J[�Ї���:��b	e�75SPBl�D�FS3��E���I	�/c�M���5���N�f�LQ��&U��:�!����*zQ�����p����VT��� Ol�R����O�B�����'�^��fӺ��z챒*�#]�K0)�g4�r��A�6 ߐ�X@�$�:��6eX�J��:�c�7�y��W�T4��A���c8�Z�C�o���Q 2�	>,\u�}����_�t4Ȃ��I�'nVo4�J�ٚ�Y18��!�E�B�Le�t8�����0��)�H��N����,�=1��{�f9�Ȏ��C���}�_��P�3��a��U��K]G�]��x�#�K1���xY2sU�z�9��4�`�"pT=e�"�gR�*?2�l'�Z�L�����G_Tqn#T$?Ҵ��5���+e-NJ�{rFM�B݁�c��!b�?�v���FK�7f���DZ�\�'ڌ�ȷupz�2������!UsWr2�-��W��M�(��Ĩ	�<���J��ֲم1�_���^�(ą
m�Q�sG�?�-p�	�~���UE��_{��3:	rkå	6x������dw�0p�Ģ�=v��xI:.�����nr�o�T��������H��w�yR�ƨF����ݖ���.^{�aFjmZځ5��t+�U�8���ՓWx8u�k��G�IȖ��cR@�Z��N�����}zb�/ܰ��Ɋ��wc���Ř��]��:��/�}����
�kyx5p.���[��!0�l�Xm�kٞ��H�(tKp
f�a������BӚ��l`������hKr�������ֽC��>p��/#I��U#��n�7R��N Th$�d�L��)��?J��5�?�f�մ-X�Ϋ���a_;���_��l����H:^���h3@4;8�pF���۷2�Tz{^�ʾt�Ѯ\�S��_��)=1O镀��{c�YS�.�'����EC�O��?��5�A7-� ��Y�H�8Sw�'Rl�Nu�N�@�W�xi�G�����$X�S	�<�0�=4�^Ӝ��^�ԍeg)PBc礫cc������z��YyNq�.��/�$�l��}���a����zVR�$�.�>�SK�Ό���U���UKR�`�����\��Y͞d�@�;#������qݟ
�O�Km#��-6�_��4��|�
�hF���|V�nr�S ���	Zۧ+�>�̕~��m'J;��Ő�a�*��PeV��a�=[�6
$W_î��i�Z浢�w8�(7
fP�
P��B+[+�m��FP8
��pd�[ح�2��z�[�*��vMl����s��iYJ�x-&]=�ؙ$J�c�`4R5G�Η&G�o8|�.n��B1�S,qx*���:��f���G{Mw�Q����� ��r�T �����F$%��L��͢�L�~M��P�4���Ir���;.˿�>M�#˶>u�J!��T*��'{l���t�@���}�[N�4 ڿyw�`�l�S�B`��pJ ����-��{�s\�:V@Ҵ`�Q8��E�Y�/�RJ2!FuA�i,�+��-_�����%K�⁫ ����<\��q��<��zܼ5�{k�L��'g�lvI^/�`6�t�L� �<~Uŕ���o�6;n�t���ʋn!iKo2��*��#�rI �/��H�����a��j�5}���D,mVd�Jʏ�Hv���'JCG֪@�ؗk��b��8��jl�)n0�IC�'�e�i��k��ԚV�^��?�:�}0�ţ��}��N�vD����
���a{]r&:>O����g��Ԟ��Q�(�7��j������|�G�[=/Q����rD�$� ڞ�kUk:��W�j9WCPr��z(��� ��r���DK�����y� ٌv��ܝD<��#�h���T���?�y��PoH�w������X�"O�]��u�p�鹾��tJL�����<�>آ�+�rUQ%F��oGj�J�Z�|9��5%��j��7���i)���!1������5��5��7D+w�������
���t�'�M{:�|��z@i�b��;�2c�Ւ�(�k'�g��������mRi-���l�����]�_`V�C9�BIJ�Kix�Y��3���~��&{�΀��7)G�9,��>�ֶ"������=� ���"�������˾&gI>��_�?@#SJ��n��~�%�����vy��ج/��DsX�� ���S�����R�Y�U+����B��RQA�����Q����Fy�|�Э�*wK����l�
E������ 6ED�AT޳�n��6o��d�ۮl����W|��n�V©���U�/����|󹔵�+Χ�E���Xyڜ�ߖ�2�����T������29ў=��O�Z;���;w�����c��=��=a4@�
NyB���K�S�d��/ګ�����GF�����Z�
�_"J*!�s�x�*��>ƿΩG	�n��_��SI���/ԫ�ɷ�wX���TOv�4���%�S9�Û1k;�	�%.�����cqk�e�M�S��l���A� �=e@h��ѝ��s
}۠q�1�َ���Liqa�-�|/J��}´�����K)N�6h�d���RM���#���K.b����I���'C��h%�D����>|;<�K�
���h�AFҔ���5�2)>���f��s�Q��`�?�
�<�����a�5��4��/B�^s���zz�I�^8�2�z�P�/^�x	1KKo�&E"тR���j/��^'���7�����+�`��&�����r��J��a�0(*���U�$�gb%u��i�3,)�E�!nG�Ji���P�#72M��V�Q}y*1��Z�I_��d |�W]��nt'��\�¶����F[��^0�|_5'5x:2�Al�H"�O�e;-ZPǀ{��~�D�� `]C��sr�|�p�vD�D|��:�����H&`�����D���|F,�M6=�v~e��Ë�� ī@ˤBYÕ1�R�~έ�AC���IE"-�f��3b�q��R�����4�
�N��.+:�,�v]6O���둋�k�2X"+[�ϋw�.M��;�t��L4���`m�Ua`_;@ H���( �~�l�o;�:���@�E������d@Y��.|�Qm�!�Os������]d�*��A��U3�8_���I�6�}S�cu�z��윓�km^�P��[~'���R�����_�썬��=�*�vH߰_Ɂ�~�@J5:o��x�P�r�Ȯn�һ�����璹�t�����#+|T��s.�a��p����
�/�b�C�����~?���ƞ۷zo�"��()���eO�֮�@>�5�r���I%�K���sN����I�%Nd��{`2� 67�t��nJ�I���+�^r��bқ؇�f�
���zEK�S�Q�b�X����*ͳa�ćӻ$̍�*�Dݰ��UZ{��� M]�%�Q~��m�,����l�h��S2��j�Q�U�W���$��g��2�L� ���0�v����J"~����p�>;?Z:?���0�l:*�_�7��dրƊ��S���-�O�A�%���.軋?��#��Ǭ~Ri)#l���(tq�*ڭr�mJ ��ӴHbC��qϫ�C�M!,n$:2�V�%�*H*�z����Ʉ M������C��K�ϐs��J�b1�Vƌfã����?y$%�w�Kb�M���&�����c��yv���$���,S�	��2�O�7S~�	Hޠbn�؏��)�'|��.���5��b�4[g(A�{�7������x�eX%ϻ�9�S��}�$�N֠N��<F�/D�k��d͋��|%��#�*�Ȝ����R[���rPXB��OJ���ף��xO+���4N��ggK4���r���T�ದ�`�|B�+Ɂ:����ئ%��
g&d�,��ާ���ėg�[���˶]�I��	�O��b�D����]�@�a��Pʏ���	��qp�<��=���&�Wvb'��h� \�x�:�V\�[$B�KJ�E�E�$���oC�BN���F������$�pK!d��{��_�c+�Il�#i���'Y�kg�T'�T|!Y�x�,��h��`N��Ω����[�?�i���i�9�����o���Q�����*�T�>�}�Plz	��(&
��|�2�dO���E���ߋ�S�ޝJO۟��M�.u�kϼ�_ؾ�'>z�+�s���G�˜�"`n��;!��%F�6��9�Kt����Ⱦ����`���E�����.�����lqg�"��58�*�Y����>�h���/d������6����ʻS�>�Y�r�e��-����҂�!���䍋ʍ�;���p�7��/dh��8�\E',,a��ţ�����4�Ȏȟ��hc��\o�޸�������(���AQGm f7���P&���j�b�KE�:5��:AV�YrMG���T��l�h?)s36By֓�Z��a��c��:�KSU'r��m���P,J1-�w<�r�=]"� �@_Fxg�����lj��'C~ְAs�}��Q��H-�����&�S�*�	���'l1PE2M��?��!�8�t)�'d,�x��4��=\<�T�(��u4^�6��*^�m%C�2��򨃇�M�y�U$�=��|��.�ǃ*M&���%�z��7,�`Yq�z��M�l�3,�@7f@)�rw�D�l�	/�T>�m�����k�9�l�Y��<�8ag�[ �>�ƌkG�q��C�G���5���d�tu9�,��l����+�ISQ�
�2�
�zG�=B�c��q�����G�m�<[���dE}}�I�g^v:���5÷�fڭ��:o�ҕh?���!I�����ȎE5Z���%�4K(/
<�F�)����b��w����9c>�����\�p�l޶È�N�GoI�����*���&{Pa&��v��Z�	4AqA�(�v|�Jq��+kϒ<�$�;@:x�u�No�|��T��>c ݻ���a����T���U�����0����9�\��Ф�k|A��z�Ý ��-�{���ő���ؚZ���)�5�E�<�Y��*!D�;���DTԠ"�/Nk��j�;�o�$���$��>.�q?C�b:�/��q��Bb���d]#+�,�,��+C�^]&ۄ0l���"߭���Ԫ�Ъjo�hɀ�[�"��'��^[2����Ʀ�yn2�!�O[�w8�e�
��^��p�$��&kQ��`�b�FJgr�-gV/g@(Y�!���`y8�>�a,,Pq	�SR��HD���;M��9_�v�6��~�y�^�b����)���+ƭ�6-u�S����5g���&��Bɨ�s��|u�s���s=���6� ���(��/�C"q����FO�#�wn�=��;�{A���;�~~��E�?;�V�O1ذ����R�T}Q��ITn�@��]����Ms�Td���w��\m��e��[�z��M74��*T ػ,C���#�0���z�Ls+���fW��[�څ\��Q3�^ͳ��P�N����*Wu�̈<}f��'MO ��������#@�`[ ������z|�~���F��R+��a�-=�Х�x��v�'6*���WM҈�3�~�:U�{W�>�`�nd(!���3�PR�C��G+~�@�b E��_��ۂ��g۔Vr�}N��K�g�{�E���ٛv��0Q�C���5�!e ���-l^u�l�����`9h4�R3*�;�
K�й�۝ ����F��b�,�;�a��PKTea"7b�$i!�T�Wk=ā�M��X���r�(?Zu�ϚO���c��x�>��N�	�r;ڦO�����V�,�PR�Ld�4�.�����7=s3��#t+O�SLf}��C"u����t�alQ��P7��γv�Z�0q��~'�Qh.�P���wMb���^a�\ r�@s�OI ����Kk��*�+�(ގz#8����pP���SE�쨧g�}��hX�$��,H�U�L�:�Ґ� ��{M��;��1��Q�kƣ��9��ֱ:(4:�(�w��4a�l[�X~(���g�f�&��4Ǧf7�F�����.�B4�i�Qіy@
곋��:�unK��ȹ����%�����Ƭ�%���G�Ɔ^K�u]nSK� `�^Ѵ�6E5���X�����~Wߞ�7����y��`M�ܳ<PL"�j.��C�ZK�j�P9�E��j��_R��0��� ���3Q9�B��45o�!�to99���z�����~A��A
R�c�z�˼���FFs�����+�UJ'�n
��=����u����)tC(�q�Z7,��F�d}`���K��c�z��!����zҡ���L��GW�٤�,� ���F�77��z�F!�+�:����l�ɜ�"���]��ٹd9C�۷� ~P�ãa�L��`�e����!���W������������L4�C��)!(K{�����ـ������)�ҕ�ąY��y�
-%:�o�'���<^�fx���<�3����ݨmB�ҳ-�����2�ɳLt0�|a9��%��2W:���9��_�!.�QN$C/&��U;�q��Ψ�5rg�x�`}FV��RM�|a#���X7�:@��	V�ѳ��Om�R�/���s�	�s�4T[-
�1s���GQ]vq����@jY�X��1��x.��;4�$��+�ڵG�'�l��NƟ��Zm@�Qb�s2�Ǩ�`'ؘ=��}7W���QRklk��R� ;��/�߷Fh��#щ����������`˓���P����s��6��Ǩw���`��P}��2��B�U��L3j%���$-�el�Żx}$F��:D�)gZ�ϭH㭹2�5�*���UjS�RU��ل����ߩVuPŪ1f57vg^��qJTp�~����@���f�!Ȣ�	��<��%�)�}"���lQ�孜�u@�UΤ5�\l�����M��7�m/�S������t���Ԡ��mO��"���j�z�	��}���:w���h�x�0�(�4 �ˢ6���W3Y82�t�d���f�ni���e�2S**��r��H��8�"v�4I*;�_���w*�b̀�����D������j>����oEUui�o���yw��O��b���MHƱ��{�x5CH���]=�����$��W�Yװ��uS�ѕ��}�L�����Q,]B��FD�Ƀg���Y�+�o���0��C��-�9ޗ ��r�)tV%���'����%P�@YE�/b-���=��N=Z��n���j(�嬶���Iˑ�2���I`.t��yq�%�7
��VMdk��.��>;f>�F��:E�&��Z�bo�^C���|�\�%t����_U}
^>��g�/8r�^"%���������Ő{�h8�I!'������?cb[�-�q��U����E�upV�l�s��kCĮ\L2N'мh��xHA�,��2��T�(��*ਲ਼��s�]ˇK�1�7�蜆	�q���▻�#��ϧK��r��+ 訓wt?C�b���ݓe���w�[��P��Z��������-��d|��'����"�r��ɳ�!z��M���)�a��Cb�D��(���Ҹ�1�o���}�g�k�g��ŝ�J~ߡQ�{� �G�����/��^����s�����A$[+�6:�~bRΣ�D�_�o@���!OF�"&k�d,��!�`L7t?Z�pm��6��L��=r�nNy��#�+�?�/CkR	)G�O�G3[j����W(�6�F@��Qq�����ּ�#/J���Qf��0 JѸ��F?�:$��5����۬����4fgp�4�^Ç��y�����@��9�ޟU#���0�M1�F���9�H�>�.M|��e#��BL�'|@�m.���E�?;�����@@f+�ʯ�@���]$s�S�����k�އ�H2�x�,���U��I?��|���ڄ�n �em����?�6�����#�02����z�i�I��mPP���?1'%y���^���_�F���Eh�N"�$7/+���EUߊi�*7Æ�WC=g&�h�������;����ѓ�`p�3��}�M��0�-�A���]>h�!"PɞU��V��@p<`�M� ���Z�M�J�]�/g���]��e�Kk�Ŭ����`��o[Жآ�ۀ��|B�e��ХНgwa�
��{�h3���RyĮ�}���ހ��?��B@����P(3rߪ>h��&��y���@`j^l���M��Wl��B��=�O�y)e��)�1�D�h@�1��9P?��w��`6��.�K�|=&g�/M���*4-3O�#G������S�U��e����r�#��g�4"b�I�j����K�.�@Ui9�|�OHL;���P���^�}�]��r3��@р�)v����$Lx�(���tL�B�ک�SA,�eg�_�(l���i�D:���I>��L��)�'(�Y��8��5��sS��^��d:9Υ�,׬�?�z�����q�(斫�JD[���VT���u!F��%n�.i��}�@���]��
Qjd,������Y��%S@S���B�%��Wl{��7i�𣏕��ǈ|��B݀⡮�.<�`��K��,�У�;.���ڑy=z|�'"�tc�,W&ʂB��(���
%���>?��Wwo����`�(��M��'x�������M;x�QgԊm_ɕ�3�gj��}�6E��{u�-_��%��V���]%�7�4=5��5%�@����+�} :���/���|i�3/�d�IV�W�V���+M�<�fw�C��{8*!;� 9,������W��Ǹ�q��D�k��`�@����M44���]�W*��l�����-K$�:���B�S�f�)�� ��'3n^6N0��Td�e d,�]N�y��&)�l�U.k"�v徹�ot���:��&����#������`�*U�<�p��bQl�]j^`�v�\��ܷ�t�Ͽ����_����hV�b.i-�B'cj��a).�b����ة���Z�O�
(#�#�<N��z��ť}�2��f�H��c6P�Y�_a� O3�2��x߇����t�u��M��p37���\�-�Ilu�>�G��rNڡ��_f`��9b�	�H�g��csnT\�����Y���DmT9P��޳=mn�xfa�7�fe_M�]8�������Mʌ�:�h��P����Zbݍ��Bɰv2k�%��23�-z�&�esb���-B��DZ2:�|�M��!e�zZ���l('[�9�����x8�d���WsLb49;t�L�"/��^�_��Uڲ�s૪U�D6�n��r���s�?y�+�;%wЉbO�ܗ����0:������:+��[��b(�>��ƹ?�?2|�U4�!�LV*�E>_��@s������/|���F�VD()��6Y�A�v�|�&����0c��2�W�Jj��6�6^�]�KR��S+a�o��*ݪ�ο�ct$/e�~M��d���^G^ʡ��1P�=\*LXCg@�#����s�f	��2�qO�# ew y&�C&�unB�I�͜OV?�9�>G�N lV�뼶�Ŋh��� �^:uG�3v�cHs��i瑓΁%�x�v�#�,���m�Vz�T���9�l�\��6׻}u�αc���	H�P�u�3�6L⫳�"�`���ho|۟��Dn��	K3(����U(�V86���*�-��M���7�)d��vG6O��k���T��G	�� nU���l�z���V>{��GH,�(�����h�9�B���>YO��+�:�<���y�Y�A>J0�MA�qX�L�,P��w)r���'F/�9����hl=����UA?,7��Vl^�l��f��}P�iۇtI.��sH�M������p96#�Q��\~��B�����w�@�~0�%k���k@��*%Y�6��غ�zE�Ew�J�l<o��ԋUg�c��a�h?y�$�pb���2Z@�����j����ܡW���?e���^q�g���߰L�H�;)-HI"�:�������YH�?f>�����!��R�~��.�o�����x4i�����_`j���)��o��HgO,|�
��7��r�L�!���q�Pp����R�M6�0l.djR�<u���rr�u}Fi��7V5I]�+�z'�=�v���=��%�,
	��Li���n�G�O{\{H�-�=�����K�� ���`�p�����J#.w/Oh�����m�ۦ�ڵ.u�k�ՉF] ��e�g�|�J�	��/o����d���a炞DdP�6����I@�o���#5V�
n��Ǫ����F�e���9е��1�+�#nX#����/��ֽŚ�Sј��y�A������`~���k����E��?/�ǨXWP��%՛�"1Hp� �bQ�}�+Y �=M9#�h��3"�
��o����$���GlV�\��=m����q��=�e�˼U*����qW-D
�adW��D���F(��i����E���a:�>;N�:kG�R��Ю�M`'�$�n�#I;M�u�,����bJ�u"�]�� 4ܱ&���b!��u�F�X����!�u#y��"�Q<����� h�@�5M�y�8y�=q[O�R42Le��)����T����*)�~��ͶXrM��#������dlX:�!��?d�Yj���S;��#�S��@�����v����8�������/CD��K���;i�F���+8%r`�	
��#^��s�B&�W��	�ҧN��K!#ۡ����$'d�A-u�Qv;%�i�M��XP��x�d�PԝJ�� �'����,����g�1͌M[�H�?,�#���+�m�����[���2o��Sl-����޳�ж�ҫS�� �z8�HJ#�L(B�D0|�(~Ec=�3?��H1jCC��ƞK���
�F��Qs���rj�QJ6q��.d%��*(t�
{�S�u'��k��ᒺ[�+���v��p2��+rM��y�M=���F�����(t��u ��R-}c�*����ƞ�=��M�J��>]&V�P�ޥ��T��������%C�ܶ��\e��	-	G�9��+�i�4Ssw�0[�<yO9�E:����cy�h��'�
~�1Ljl��bp��PE�r��C緍(��:PA�Ի�8���u��Z�gu���ܤ���z%( <�u�B4G2˰:BW@U@���r�f�C�S�fE��d�RH�G�g,�80r谇�� �NG1 5�ut|�mӞK�O|gQ!���..�n^��CO�����q������>�����H�]��#���N`v]�Ha��j�p�h����+�m�����B���\�S|l�\>>N��pJ�����W��`)���&���T2 i���#u��2{tsq� ȩ���v�����tu�J��j&�sv�y��vȒ��M��,��/��ސX��PN��%�ԃh�L��OU}O���w�#|Xڈ~��9��^>��t�����	EDOJ�9��|�k�V�YAAJ�O�-^m@@F����ya�4.=$�e)�,^�p=�@�Qu�p����6|�t�'�@�nt����Z�}nvߣ��.�	H1��m�u�Liv�"M���u���?}ޅ���+�h3��W���$��IzO�M�:�$��O�	8Ͱܢ�,�;��~I��3�j��݋ �\���Y\�I+Ω���^{ �멂W���g���4,�8��: F@"��0�Ja���&v\�1"2�W�/�����C��(����w`�uK���������W�����5>��ӿE)��A��Fi�P��������ʥ�Á)�	/�b��5��ÛffSS"���m,��/���MT���^2wv+���6QL?o�F��k�xR��U\�'��c8�f��C���T�i����e�z����F��9�);$���H|�{�e ���'��:�m��H�Ip4�򮟾�Pbv�?�V9>%R�'ƭ",\��J�3��@�q��D�-l<�V���✶~y���H
�7�Y[΁P���Bo������	��`�L���\ÌM|��
.���}�M�gtX1~\�8���H����C��\�&�W���
�TD�K鶎14�U��0N�Θ����O��� :�5��U�0�&=�l���4�y&u�R�K�8�x�
R �ޓ:�U9��R��>��x�ؓ��,׎�UG�Jx�?�5ׄ��{��}�`��k�y�ב�}"�&sJ��~��gۓW�a���W��!ۡ��0#�s�:Y�9J<�у\�>a^椝�R����]�1��:6��6��U��b=���mp=L):j1�{b`N����Aϔ���0.�BǠ� <�4h�"��Y���D�٠2��8���� *�ϔA����3�By�����.	�㗏�]�36k㽦6X���e$0���=mJP^Յ�IcM�����ls�c�J3(�՝��;!�<��~��. ~�� �̜�{%%qG��4�N���T�
8�v�"B�VfwLi���<�F������`�D5��x�0(
~K�q��u/C��C��Nh@o9����L����
,`%s��p;$�����T�ݕ���9�y�x�p���	C2%e�3�l�&x���ڿ��T\_�m���!l��X�� �`/���
>��p��}��I���߫�w��ۘ_!E<�z����Éy�I0:����O����2����Q�b�@�����5w�_~�B�e�*A*���%B��p����4k��Je��F�b�8�v�l�r�;�5����+Ӹ��z�W��υ]2�=�D¶rw��p��UX%���`�d���#�-<�w`�zca/���)U�9p:�2����V���l
��*��"$Y|O��t��4�;A���9?T�1�?�&:�X]�,̴�.w����v���g^ɚ��n�b��]�������	�4X�n�11��4�i5�T��s!~�=(_�2Ň�Ja/iR�|�����l��\P�AJ�����Q��0����=W��w$0d�)GwP�<��q9
4CBKzǶ����ur��0�h�>����:���<�h�&�d�s�u�Ԅ�����V�����V�bA�Ȩ�il4�e�]��Gʹ� + �g�NMI�Za���Z��w)C�O����� :����?i�OCi��G�^�+�T�s�����0�"��Hn0l���3���-PYcc���!uɏ��x	�2���V������=�|�SF`1�05�N.as9��Z�Sz��3��^Q�W0��e89�k;����ѷ��"WKgDՁ(��8�\On"~�(�[
!iG�{�y&o�`�����r��,1su��GM�,��x�GYK<���&���E�.p�Q����),�?ە��l���RIjF�OSx&��;���`&��L�E��;�VՐ��� �� ����g!.;a�]6�m&�l��"=
4�ǡ\=�H�\��P�9��v�A)�q7h�6_�QF��:��_`������Lj�D��`ᑂ��7����U�Y��Ob�d�k�DW+�+90���UQ���f_�rxF빚�O^�'��|�1��Ǝ�K���f��p���m�2��<)�������ol�ɴ�\h {����6�}0yҟ�������+�$ךD9%�M߭-��U2Au־�|�v~�O	@�*�٪����F�F�<*�!uވ?�x��(�����:�04'^f���>ᖉ9i�5{� �Mb"�q����.&�jG�m�ȷ�>`��?f������d��#ֽ��R�袪U^Q{#)�5J�'W����T=�u�lW��"����� �J��"v�WgNrK�"����C��9d�S�U,(�R���� �l��ø�]c@�wwh:�F.
�	=0�|�{3Y&OeT�ϐz�a-'~	Y��Io����M��)(5izƋY�~�kK����n��ɧ{�?�&�q�IU���CB'T`����9����X��k�XJ`���P��q�~���^f��.(҂��d���Ȟ(x"G�������h�H��ĉ�Q�)�A�sb�RyLۤ�z�&���D��nA
���蒳@uO�X��U
5j2��.1���0�1�%�AfUꫂ�4&I^�H��VИ��r�t�& hMpNF�9[���A���]V4�S���3HJ�1�q�sg����n��h��PA�H�)���Z�T&�JL�).���D~�?O���5.L����eOX��>�FGa~Ȣ�|���=DG��Ce����*��nS����J���¨�9�*�$NmfK�4,�-"�:����Ǚ,CD�u���3_O�f��@�A���&��<�x�dH����}�W�+M��l_(�Z~��8W�~hFq�Wn4G��V
���ֺ��~�<�W��<)L;�Y���\{�5����k���e�|���p����؁Hg+�M�aǼx��z^:*X#�!ù������k�wh�Q�Z�$Ϝ�/��Ƨfwh��h�V��7	xP�Ud���_K��#om+��f��3,M/�u�L�W6�:Ut�O白#��.cގ�d.r�� y�eι�fbR��P_s��}��nzQ̨������\P�t�Jq�5g�3k~E�_�ֹ�3����E�H0��2:b��%�_��ӌ	}���Fv�x��}����﫼h�@���~g&@�u���`PK��QS;��\y�-~5 C3	j�D���Z��MI��Rh:G�};�{�O�aJ�\&�M��+3�g���,g]}$T�k��.tu/����h≢���F���"�V��[.���25gS38Q ȐF��8���"n0�c�A�ch��Dĥz�Y�<��έ���A�dm�2��V��[D~�ɐ�����À����5�g�aK�/80�CUW������u#C_�k�9�`�+1��
�t�Пq]Zvȉ9��o?���m�n�_���8%��!;Jդr�ӠM��xa���j7 D�H-YR�~O�m���o�Ch�f�MO�
}�ٱ��Oܥ�77�%
pzwc�\g{�:xT���h�PY�!����@���
��.��S9��Aդ)������4q�)2k���_�_�tZ�k��G6�0���i(!�RU��HQ�ȏZd��v�@��H��^�$�m���BI}�c� ��-��J�R��H�5�������X��Kxn�-��%�����)�r4�<_�0����fE��|쵲C"�n���J��5�	DNi�G���CQ�)lu��w���(O������8T�a���F`������٨Ir�: �q����Wé;:c�<ދ�K4�\�7��"\Ym~�tC�3�(��%o�4;¿|<��먻�nC�1yn�[|}Q�;L
Y㙿��Q�Ae�d{�c�R�@e��t��<0 :R��oRgh���`�C+;�'�mw��<��/��N����>��G6r����5/.)2-�$(�i����6�Cu����1r`�e*\��Lp3�bz�V��-�Ӣ�������ժ���*@E�7��M���G�^�� C3B�Ј��G� s)MU�Q'r""��vp֎���,h���ō��H׷NK�^�	���:��5�J�8>�t�wB���)���!�ڌ1R����C�Aj�Щ���iE�8�բ���'�'���8R��_�zֱ�C�G$��!�i%`�����y�����Ƕ�����/��[���$B�c-x�3�2�t7Eo����6�;y\�*W�������Ӻ�%ƹ�W��]�&Uz�����ʉeq'��O�	/7�V��	X�E��+ऱO���D���{�~DBs^_��Xߐ�8�I^�"7is:'��#��:��zj468%���]}���;�1�sl��i�G�dϯ�^A�㊮�_YT:���3?[�(�G#i]�i߲��]���/?��Ww?-F%���]2�i��0�0�-�1L�|��h�5�KfWB8���28�t1��S���bV��*fز ���r�E�t=�]GD�T>�L���_o�B���<[U���[����}~�@P5��	^�L���`���UE8n�-�(�k��O��M�PϤ��4�}[ꐌ�����f�8վ���7��)~n�p�;F6�-_ߜ��T�V�l�4/����M� �ZDo�_qc��Vo@�X�r����w�f���	�VH'<~N�n�,9@�]4� �"�2�1O�m��T>�?./ #���UE�T�TVE�K�L��1G��^��&���&p� -	n����7�ې~��b��`����.j��1��=����	T!�"%��445f���-�cGRd�n�"zG�$�Z��v�$�$��ml�~ ;c��>Y>M�x�0���	��-����a���ͤ�R�w�.
|쌹���1+n8�s�i���XOc]���7�
�:�6%5e+.NwR��ɥ����Y�72�^��=\7���Xs�m��ɩ� ��*�Q��&��}��e�UV��9�3���U�&����r�Q��?:c���~�dF)�B����W-��LQā$#$9�Kr��j��z�Y���1�p���x��vI�@��s��z.�gR�W"� ��]�N<����ÂKJ�Z�q�Ѣ�oگ�X]y��d(��c��6��y.�S"��d���#A"�e�V/ߏ��&��C{�Z�2!�#(Ɇ>�R��&<$'fH�ݡ���aGS/"j�����b���𶷞�\f�����R������9���Z��3�C!�ٜ�JK���_�D�11��_����d�bE�r�����T;(?9���E�uEJ}~�Eڇ܃{��5�;�\N2�k���-�P�J�	�1�14�|I�S���$Z������i
��ژ/�k\Ю[k�F�&kL>�x�u��b����^��G�Zu��g꽠�A��
׆�|��-�걻`�	]μ��:+�_	�E���iv�L�diu�$�N/ߋ?X����) �����z"�!L��j��4F��]�ڃ��)�ZI���`�Y����Ϊ�&ӂA��8
=*��!�#��?����������'��S�*֒j<�e4g��ɠ��7�h�>��E�'}	�c^L.4d�(�|��*�װ?��wF�eL/BS�N�U�L��lP���1���`0�W�e��pLU �x��Qd��TT��E.i�P�����n����A�R�����"l�G��s�EL@��nC��&чN�7~�0�Gd��k\"ٞI{��`����Ce�K�a*_�L�-I�Ɲ	&�Y,�yEK�� ����HR�t㉕�F�, �Оqҕ������s6�U�Z���u�H��	&�h����ˆ-F�X��&̋b��־�i៳׉�������4�W�cT�R�l��ͺ<C������C\�d?���i��QL�Z�	�1 bµa^X�ct{)�6&g1��np_�}&�_#���܁��l]�����Ղ��5�����8K�82�6��j�uc�Q��O� ��7��4��U�1F%Kii�V��/�i2����>e�/����A�JH��Z�x�ٶ�?����l�]x��v}+]�H���^���J�8^l���d��-�D��U9f��q�Uւ>
`�����Ū�:y?�x�t� T�jG�W�����T�,���c~ZɅ�E[����9���$]��� �|�ܣh���yQ� �&X����U���W���R�-ݨ��eE��L�M�ОE��ύ�S-�?���6GB�rNd���!�<���ؿ�r�8���mF;\��WP����lI>�ˆ.i�D���J.A��4QL��|������`��7��(�27׌{n_��z���G ;�S�<�+ߟF7��#f�x[�x~�Z��)����+W��� ���5Z.�4�RD-��y��n���o�t��@���/Uy'dr� �pl<��9�TXPmRM�v띖�������#s>�01�L�|p�cK5 9B��KnmK��dx���P`��1��Z�VMD+4���n��-�񑔘��_�b����7��Z�Z�N`]�C���n7��1��\�pn�|>���Vo��5��Ǉ���;z��\<�Ra�8�������ź�;ZPt�n2M�oV��JT9!Ѳ_���t֩��%�Y����ΖP��e-�^�=��؜KҒ���;a�a���
��-�:X�I.k/TU����e쐚��m�9�[�HdL��2(��� B�ā���#N��pf4KF�k�xL�4�O��τ������+��:�Qc�wkW�J�6�(�"L�q"$�RV��P��d�ԡˮ;�V��P�JZJK��e�`j���AfS��0[A����h�2-�[=c�l�ZS'�<M�A�/ �'��ed�������
�|������MV��-�
W�+%�X�m�?��j��T���#;��r�N���<�xR�#d��J�H�F���a![d�QD\S�?VMw�T���I�.���t�_���&�xo��a���v��e�$����=Ĝ���]ʫ^��ҳ�� �j2#�u�lU�*����I����)R�E��zj)�ۆc��,p�_@澴L�{�n���&�&��NA���J��,O�2)h����q�n��yef�õ ��E����
9t�s�e�e�C�E�HLLg��sئ�D~����5�^oy\_�γҫ}n�Y�{ۢ��.� ҇3i,R)n�RbO���@��p��/%xFEQT0�w��V[F��.�LP�9?o�JOju�xYv�-�%�e��������'���b)���)�ηP�~O]�e
���襩�?3�`�O�^E5��Ծ�jp4��RF�c���� <�	�:ڞQ+0q@�Δu\�-8-qü���/+j��K�Ӳ%��#ޱ^�a�����
{ceO斗�l� ~9�`�_��#F#u�R-P���� �~U63�8_s�]%��R5bZ�۷v���y`k�1��|��=&��QFN��R���MҒ�Π�Ap<vdrr�7Z�[��F�������ۺe�R�O%��x`Ip"
<yf�G�&���*��A�J�y{����x��3%,�ɍ�@�YM�6E0|�!Cc�@�i��gb��>NҠ�8%����-#���$(���-�8s�0�<�L�R���M���g�S�+=�E�TC����*W���Њ���C��e��Q�5ڶ�_<l�*@���i� �����d��EJ���lkQ7#�mɄ�  �G�����/!^���F3�T��8��}�4��Kǻ;�( �n"&�B�Ǡ���������e�2c�U��3�o�`�9���_i�u;��)�u�ͿZ�m43y�c6��o!-L�V�F3�9zZ����u`Qb��u���E.}�6�ю ��R�<#е�����5d��;灨�u�g��k���m~�R�Cu�VxP���ـ����N`[���]% �'�2�*.2j5�l����+;U��ȠE���� ��ƾ'�j��ɡ|a!+no�iD��B�{��[�p�c��{�s�U����=
"q��e� Uf�j��K*3��px8��E�$X����u�#�J�g�31�e�~�{��.����k�x��Ә^;p�n{�vz�ȅl�W
6�ёn\y��]�$74_H�Ӳ/#b���.�D/[�]I[�M�m�SzY��i@7:�я�s��s�e2&�AI�����RD����N��-��;�qj�zX�61�bw"�I8Z�g�>��:wnI�7kyfACz�uª,�L�~�h9���亸�r|�4xȒ,d\�gl/N�����G3$9A��cw�t�FW)y_\>twNo�Q}Rd'R�Vc�� GX����fr��t�zCMQ���	����lTȸ�	ڂW�da��H���+9�<E�?�/�b����ي��9�۽���	��B|�}95!��P^�=�Z�G�޾@Ri��P[]�j��,�D�_8~��'����o�^��j�H���H�F�\V6��/W�uk��j�&Yd�8��~A�<�cM�`���.#H{m8d�
��d*l^���X/�<�t����ϩ{�72_.E8�P�f��Kl��WȜ��ryyۭȹ=�L}s����i���.�B�-��Jz��@�9l��i�ⱇ�Y
8�?��	�m���?UPd���S�k>Rr��y�Om�׋H ��S�J?;�<s*�U	������-���w̼[�u��O�E"��`;~���]��`����M?j�x8 +]&�tt.��%Ls���&�$��̃g��&X���+��~,H�����C����`c��}!.0�O~�%�KR/Q5�Q��a>�	Lm=�V�խ^2�铁"��1���� �`
�&�[��T�W�aTɲR���Z��=�\!�-�l����{bg)1[�K��zD�g+!�w�$��
e,�~n��O2� �v�$m��Q��U��K�E �T5@wJ�Y���\b�3�S���o�k��z�@�#)������T�ry1?5��`�vxf
��%�@��b��@�������ө�[��*���_�)f�>\��a�|_�������)-���"6-�4��t�aY�T׉
J����Uи�7��y����g����qΐ��d2�4�!�����z
�3Ov%7�HE�&.���-�o�F�Z�>���5�E���PoS���=��d ���U�O��r�14O���d��n��x��t�d:��MY.���l <����mtmir\����#����
�)ڧ�?�X٤?����b��e��~���?�q�l|�eh��@@��R�D��R�&\s��[���bo)�9U���s9A"�,���W��6)��}��uoWXY��������C�� C�*]����G�L�{�5��a�A��t���\���5��x.�zd����y��}��N|Yos2Sd�'���Ý�+�B�W���߰��Ju��?�k:��'���#l^�Y�F��Kkfվ4�էZb���!^8Q�����⾨��3e=u�-�'np�N��\^�D5���i��3�:Gt�es#��p�����2k�O	 �b�r9Nz���8��� ��O>䆿� ��@�4-�]C;�]]+{#u�>�*��R�^3O��d8yWo]�~<S�;���ˠI��cC�Gjxzd�V��kU��&��J҈+�Ip0�6�s�i�Fg�2)y�	_	@��Y���0�/�ț�� b;l�i�S
䵩��X｣;��q�9���2���׬�C��O.]���#�����ބ̥�&���}{3K�h�ֲUl�����!:^{\v��*�#��t��ϖ���ū�v�Z���!�1oY/�Tb��������-�#��!��Β/y��p��dp�s4�=3�;�+�!�(�hé�l�AyU�?D�Ŷ�����=0-����ڥ|.��q0�u_Y��!�� �	P�<������
"�SyӶ�		��v������KȎ�^f9Ui*��v߮��M���l��)�̤�-��MЉQ �d�za�nm����"�+�h�&m��,FC|���$Lp�)��#[�h�S)�)+�����!#��/V �����B����ˀW�Qsa�8vp8xu�
��j=�+'�A{�utO*�.��O/n�i}���Z?�j������=sZ�� �<� o�t�`ɞTJ��;"��$�i]���w4���R���
s�������^7Ú�N�Z|���8�u�h�#{(��i��5�Sk��`vc�\�%�B}�k�N�MJ�np�ɏXf05]�𷇩(��@,X�'��˶l����� ��
dEʢ s`I���&qP�ǥ�<O�7�h\�����:��<�4�ݠ�f9@MS8��𿶦��N�b!�����iV�¿%c�h$9�C��X�wt���ў��^�ֈc�^��I���Ü���!�u�5���p�ݏͰ��	T�=�`M»|�bp%6�(����[��M\�ϒ���[�~sH:M��r��d����OF�LvR{�ȡ���C+�>Ad՚%�A+�g8�/G��g�����/��L�%Ԇw2�`Ub���ڊ��g�Gָ��e��} Q��$	�o�U�PU�A �j��� s�p�ˈ�&'��}{�X�1��O>���1�)+�J"73�
{�Yl=�jA��z&��w˶�"չ�M��j�Q��/��y?ijo���V�[�d�̌���C�l�</��UH!��[�|.���~@W]q��Xܯl7^H)ɬ�.��@n:NRw�ȵ��-��'�	 �7V���F1B�������K�N����,�R�0B.w��XB�B~j�q�,a�c.��H�%�sA0WI̓���
�m)XH�/?��9��.Rd��JZ�`��RA��z#ʹ:_��"<�o�X8;Δ��J������OS_�h��D�Ќfӻ懅��L�V,�Ƃ��w���V��o�pŉ�����-�6 �e�,�,l���ҧZ́2�AA��x6��J���W��Py�<f,�.؇�=㋟Vم��PXX�!�����ڃ���:�i=���6�(�$��rJW9��7�
F�`B��r�,=X��%-/-s^"�I_顬�sW��V���.��D)��3��� ���)�9���'�(ʐF�;�=G��_YM��uҷ�,4êǍn]^p�"�R� �f6=��"�]���I��m�v��%�d�b�$&�2�Nu1�3����bU����������M��[�x�1Ɂ�9 *����qn����[3�ī���v�$i-�@䞢Z	'��S�C��`��X��~ώ�w%�������\���*��.�l�n.��^k
)��s�a�W<B�٪Fh���g֬�ϓjMt��l���$�6�~�ں�ը�O�a���Fv�"��)��6�<�/z�X�d���t�:�<G�&sP�}8@^	NL�:6�)N��F6�D�;�b�����j��E��W�!{ız�]�7���KD���b!�+��
���b1E���F��yQ�/�{�� 0}?�B�8��{O�5,�Ȣ���@�^��:�\�*}{��]��h��=ϦzY�zU30OF6�B0G��s�8	=�nKJ�=ו��h��t��IH,w�F���b{%�/������yG|�A:�v����]�}�Du��p	�8>�[�K�MR���b�� �(<��Y�*� W����V�e}�G�x4���Mf����}"�z~Q��-�0{�d�ySȭ؇��veÐ�v�,@�S[s^}����a�U9:)F:[[��`MV��N���n�SN<Po����2P��� �ڞS(q��<Š�eњA�D5�S���DEk�wy��V�*x��'w^���N7�qڗh�%��Y,袀�Ű��
�����d���Т���m�Í��w������%�c��p�	��|mTGP�e��ܔ(*�����i9&�q˳��.Gj
�W+CVv=��yx�@\���=kge��8���I�A%c*����ʥvg�Z�Y���7�&v�^�k<ә����
f4��/�I.���^x�0ۗ|����o��_���� �Va+� �j7��X�
2�I�u�X�TDM�����c�9����5��Dz�_�w����)j��4��ZÇ��i_M��^��l� sA:�Dn|�LR���I"r�~�����+�K/�f	���1���jy��V �Ҿ��O@�lm
�>���6��sD7���GeF��	��at�)�p�.h��-4�O�n�T
(�#Afo�dx)f�t��κ�Fl��؁�m�$�[��dt���	�鄊w�1�q~���=�W�ְI�R����If�M�.�\kn��^�q<��UVE���$�DF0�Ey%6d� `�m
c�T���ޑ'��Pj-/�����:E�#�'�Ë�����M!В�"�,�u�3f-��'�W#@�g���ʾߤ��%~�.�����<F޺���I�
~	M9�p�\�vhg_��Ε1��.#��:n���fv��0�BV�(C�����.��/�Mh��B���1�e�v�a{U}�T��΅à�>���{�ƫvKt3o���3lqj��� {n,����^!O7�ޙ;���Kt��JUo�I��=(j`g�!��2�&߷��O;N
*j��V����le�!pn��h�:�Ұ���<�2d�����"��/J;p��U���{��,�T��	ȏ�
�p�/��П���67�@�8�v?Iu�E�P��qGx��,���-	Rw��&����qZ�(W��oV0>g�� ]����,��	�U��1�U||z��ު ��z�A�X�`�;�1 4{�u�� ��kc�_zmm���^�_���fAj����)����C&6ᶞ@����[fթ�H�o��sK!@z�J��jMY=<�&I�ܩ6O�%I��hTW�.w&�m{q���;��EcX< K=I�슣���1�!�ٜ�y\�j�$UV��JՋ_U[׳��/��V)�*�qѭ�f��C�M����Pl�$�NP��Թ��P��K��B~?����
�8�I�$��Ӭ6W�þ�:)G����~����A���P� ����i���3�Y.1(��z�o@��f��6*~���2K_����q&Q�[U7�>qN�3(?kgL�v���N�Ib�0����/��+<��E���Ҹ|���!8mi���sM8���n�����Al^���:��M�c����?��I���j�ee
Ax�n���΀���$Aw�\M�xԗ�|�?������Ï��"��Ȅ��֠Lx3s�SƯ��G��B��:���A~�j���K�G�NH7;IE,Y��n� �3����'F3�'�[�u�#1h��0�A^��7\g!!D������I�e�)#0è��%�ցϵ)����7���30�N`Zx�#�Ob׼�Xk�㖇��c�Ms�����'�F���#�fH����Z\L��4�JjW.L��W�N��1�R�n>������E��CJ������E��B��M�͡���3��o���
�8V��xe���}#ؙ���f�z����<`J��}�r�T����� �`�n�sQ�+b; �{��a��;\r(�^� ��Z��-e������f��Jc�5��{������{���c�F��gQ������)�z�,$vIY���P�|�P�>pf�Guύ�z]�K�b��s��4�I�� +�Z��\�b�E܃��1S@�V��֞P5�y�)]G�H�E�?|��.^�����}��&x��R%�� k��7�[��UeJf�/#c��KjA��-#D+��)��u��^�޾�jZT"���2�!�/�T߾g���;i�sU�5���m�/^�p�mG��-��W�x�H�%H24��a����J1���E�: (�p2`�(�����8�yP!^�u髏9�zVU�e�/t�Fy�Y��~)�K!cT����`?y�XP'c�e��$u�"!�X��rtI�B[�ȗ�,r�{��m}����g���$}`�#�Jq����/Yo>;�sD_��u@�=u_��@3��g>]�t�A@��˖#�d����T�?د��;���`��Tݣ6K"%ٝ�B|<0\�9��(�m؄</�'	���?�����U-�p~u�f�՚#jl&�Yq��E��b�q�C������Hs1`i������^�=���b"e<Ʃ�:�����s�E ��S�7���C�yٴ�|�Y����')��X��WY]���	�H<f~H�NŊuea�\������`��S��27���������w�����|<Ȍ�'k��0��vj���q��X�Wt��?�o����ݽ��ߪ3X��BO�|qq���$@� t@[��ԃ� pÅ'�A2��]��=U��GCƔ@s;;9&�����x{SC8�JZ�-Vq������;�ˍ�L��"�t�=t�;��.�^���T]἖T�B�7C&	������u���׭g�Bm�x4�f����b�x䣠�\$^��yU�Uʸ��)bH�6��@��~g	r��w����;4��tH��=Bs�a?=�1!�3�//��Hg�N�:EQ$�p�ZZky�/x-���~o�[�S3 ����Ƅ�Y�X�'��oa��`�T����4�`xEX� �S�2�9���";�eZ����h]�E�}�FD�8��{�P��^�ـR����zBy����HӟV��Z�*��;u[Qe��7O�S���_�X����h��G�������#�w�r���Z�P�/�a���{�;��5����	�^X�ܦ�xM>F���S�/�42b1~$��CY�����j1��m��8S���j ��P��ߵ��=�T��vQ��-��J�κ2fZP�֭yt�c2�������J BƄD("���CT_@\W�]�����p*�q���x����%�"x�OI�}�|Ŕ����M��?%�o�p�#����|��HNvx_�5H�;~'%��u��h�ǁ�4�����o��C� �z������5.�G�E)|����:2%�}W�������[o��g�Y܋;�%�{��
,�{�<���y�81|x*/AW�m���~� �}�P���`��W������)�I�_%:���&RTs�o�Z'wb�3�.�jϋt,W?kR��' B��5���d����6���+�f��!��;�7�;1F����y���;�j&7�Qz�O	����}��T��D���9�	��Y��ܕoM+�
����yGc�w(�g��T30�W�|u �0ۈ38� �!�V�ԟ�/x��T^���QU����$��9�P4�f�8F�Yr��Jze�{Ԉ���3��V.v�j��7�����oN�����1�|K���r���	���p�|Y3	=�ӤjO1K���c>�h�:�q�Ĉ���K"��U�[��W�k5�e��y�ux��ꋿ�#u�����q����&��Ӄ�Jq6����R��X�����q�t<E)���M����/�d�g]�_�CĽ��i��3)?~Tĺ��ˀ��9	1�Ƕ��D��E_	b�86�����j}s�p�2���)��J|N�x5�ĵn6bD$@����Q�ɱ �cp����"��	ƥ�t.{�(oV�]c�(�������+�����zh��2">``��!��b��LaX��ciH|�6h��c-��s�5�M+��)��ł�v��\���k�_�x}��W�P�^ï��̕3D����F��-�ם�� t�y1��Z��Q�3^��
K�{1uG^S� G*s��pT����%���~��zz�Ih�βҼ|� ��c�>x�q��7�UN�E/j�$/_C���2A��(���	r�(:*���ico�m���E�gl�nl���<��{�D�Eo-T���(�x�r��хU�,���O(ُUl���������o��%,5�U�g ����BϮ�5ܡ�����f(��Ԟ=�۴��ǲb��p�����2�|$����fz��B1߀�MW����z��E�-�녥K>s�g�Hv�ui ��T�Ve�x��@h(ܸ���ִ{�O�I+(���Zg�AP�C?��Iނ�oK�!R���?@�X�i4��n���"+4��͖g�$;�ܱ�[�ُ X�]��o��*E�<Ms��,�j͒���W�>4�<[A��W����&�v�I�ϓ��W(;cƍa5(���Z�m��������&QN��V�-4\*�N��`!��r\Z'2�j�����̢(+���|��&��r��uQ���N�=���%�7nـ����\���{2Hd�\r�H��zf������8����w!��Ӆdv�B�q%���*X�^W%����W�C��uQ�>ψ�L�s2[�����A�<5��M	�����x��_ϛl�\�ܫJ���������:��,�	A�s�}~.�`���t]�� �ݍ`��y�V�.�{gDJ�<,+�p"�٣��\3���Y�׺��&�������ܭ�� ���âỚ�,��s~nzJ��ұ��>'�l�����d>ϼ�����[,@��ë3�$��(��m]S���([�\�z:,�KZ@�o�,�ük�'c�1�����/`�b.��(xLrޥ�Xi��?�m8���r���ys)�>��hN3���/��L$�N&�%�1��U�3͐L� �=�.�1���8?1�xS[��&L^���ّN�Bڙ+��;���y^�n�d�3��z��
>��R�2}oB��/�:���'?�4�j*Pm(^tnq��\���{�J�nP�Ѐ5iL��@m��>M��o�ĭb�5]�K~��]��o�h�5��^C���> �wz�Nר�#R�jQ�,�������3)��.��˓l�!,���ҥ�"��F'`��x����7 D\�mQ�(1^�AL�|q����ou�f�`U�2C���J���0��Z��^� ��ty
Ի`�Ä#���!HMMb�L`sW}�.��_#D���4}��
� �W��<�uf���͡"X����\㥁����\m��<�A�������T�!ڼ ��Wު�Y`���I����U�z{H;�cG Q�2��@�p�rnd�ڎ����I�84}��	*P���h�wߩxX"m�	��fW�b�O�cw�N�+:E��乍�*�v>���#i�9��M�,C���`�H�e�[w�����Pdv��^���k�Ә�m���� �e�F uAGAr^J~�r���)Q�Fi,��iǞ �R��=IB��(���DT#_ �sNĞ�qQ4i͸9�}�$.-�4?@Q�/8��7�ױ�������-��{c�u�8%����� B0.�H����1
ZF���[!�������&�}CB�|�J��h���(��&�s��	����&*�L����X�0�V�e��o��=���i�hY������s������vo�IS�G�����-�X�f
�T�W���f(��z�H��n�w�\V_f��4�Ψ�q/\�7���t���Z�����f�[�\����[Yx[�l��$�Wz>N+!u"@L����[�{xM�&�bk�:�o~��G�Pd�T��|Kr2�t�*4����OXG8��%�i����@��3���W�@׷�
j-7�7�i�YՇ��."�°~��\V����Ndc�U��:��Qe�"�7�>��᱋zVq<}��C*41�+�����*�l�I�#_z3�!����\�6�tL2X�zv�ك*���b���Jc泰�2����|�A���z��5&-";�C��4���d���7_v���f��� T������/	3����(��Ѹ��/� &�=���Lآ�M���r��!1��-�f���J��2/� l'n�D�RP�f�����]�O��z[((��]���|��ī�~�%2�����̪��4 "�,����"����F�b��r($��~��Z(�� �YӔZ���SǶ�9uH²;rӵ1;��[��Te�[s�&|��j~��A�$sr���2IP��R�����M�ǀZ�->h�Q���L��~����sR�Z�#t�`��-2'UB���4rn8�f}Xww�ڒ)�04�@�3�hZ"�����/MPֆ,�|G.x��W��1qb^�|(?<���m (��sK+9Ǻ���t�vׂ
�F��&�������Qa#��+�\���1\�d�����阜b>�w#����~Сvݿ�䐡�����գ��^C��Eȗeذ+a��m6/�'�����tPq��^z�<cGQ���e>�X@�i��|���� �~�6a�������"^K�M�D��.�}>�+�$8˵��KHR�~|߮��>vӁ�8@́�%k{��W�2܎�/���e��*6��,+RR���u���<\������Ŵ�H2���T��%��1�2��G�c��$�9��` �TH2�8�ZR�����&_0K!Zς�$��|9�������#d����r��.V�F,~�!�d7��j�� �4�S7B伶�N&�&G�k�W��%��'���߼��%��k~�s���h9��eJ��ߞ��� �h�3��`�-�ToS��@�E����<6D�,���:rz�5ӧuӧ^/��4[[�@���K9��-�q�ɵ��KA�|�8s,*f���]��hr�g�K�5;�ʖ���:�5�noP�L� 
5|��Ub\/�ߌ����U4�4��Pl����pg��C��W�?�x��� 9�_������b����u{K�/u�^�8��D��$p��OG�{�g������C�CLAe 0�?n>[��x�^a��v�[_`�_rq�	�&=�[J'��O�� ~��aM�AE�x����g8�6�53q��Wi�H�٠������&�43�
��W�hѡ3�y:{y����|�f%�!���p8�a�YW��қP�G�)�$��Y���v3��D�V�ݐr�+��<P�7)���_���1�h�tS+h-��@m��.c-���!�6��r������t$�^��ͳv�w���ۼ2Zw杺c�\��]��]d{�#����_�%P�!�dU�RY�!��^���S��	��ڠ+�g�F�w���w�6��u-�gj��1sϏ1�5*`�E�eV֙�$@HC٣tiMl0ʩ��|������7�C�S�^�D��X:�;��MI��cC8����Ki-`�fh>���ʯI�VL|	�%'�G�?>F �-�6�H~���y�2��C�p���H6�e�;��'l���qŐ�7�6�o>����)�OE���N�p��D&��}�X�� &R����+T��e,�	�z��R6�k�x'b�����=���ܴsF���I1��`�,�w�R�]���Ƒ����ÚO��z�����[}�P<��}�6|�T*`�:��/�m��翵��R`�%3�I�d�YF����gg�d1����E�<I��Wւ S�r��x�)(��Ƕ.��?D�옔���W��!3������5�pY ��T������/k9tϏV�|q�n�c��t�h�|rF�F���h@�jB���ta!��� �E���5*��F��a���^ܰ^ͮ�h�Ob�{���k���s�P�|ՀƠ�uv�$��GH�:�V֏��;�-�vq�̒��_��tm��j_쎐&�EG�*gm��I�a�J�亿�ن�k��'��Mi7*���A��u%Te��=��-=����şa�Y�O�`�e��K�ջ�	���g 3͹B��i�S��5Z�ED+j�|������9c���9f���v���'�e����*�b*��ڼ��	X���TKϻ@ög�D3t��6
��yi�xfg:z�{��JT�Q�K˫�ȸ�g�������*����bڤ�&#Mk��Sc>����z��Wد?�f�F�.���aN��m��:�{t�^��%�/��]�ϙcPp=8E����c��x��I�=��5�������|�pC�''(r��y�T��0�t�Aٳ Ɇ�g�F�{�i��u����<�}�ϟ�����v4�[����
P���zL؏htp-}�Kg@/�b7GaۂG۟Q�/f����W�~l���$��닢q=�R* S���)g<��1Y�\U�P[���5W�]a���2`�����[;�mɱl/���`	�d��sjF���	t�Bg���WFQ�Pڳ>2���J�~��}0�w§�1�#��t��ݾ�A/g6���>�{;��ҢO��3�(Ѭ�^��z��J�6�ď�55��3�7��>��H��#һ7���őÉs6�OaxG=ڗ&T7Q���븮����j�M����F�楛�n����F��i1X�<7Мؘ�����T���]���&����VF���h����K pNyw�)�k2���Ҋ~+��qg:(z��{�=$Tj��-�F�*�/��f@����	Č���}���
�E�ó
����DY q�}�)AB�K���Q�G��\צ~�ӹn9,�w�h3�������a�Z������o��?��y���t�JsB��E��?/��٧E���K��D~'f��P���9��֣s�3�-/�	�F����e�ߵ�h��Əf�d��nx�:S`ŅO펅��*'��Jk{+J )^�ڎ,Gظj�{J�6�A�6~��12
�{��.ڊ�zB�q�c��EtY9ѻߑ� 4�4����% �mD��~J6X��r�$���y ך�)����`s�ť�]�J(�iR!,Y@��Qѩr0�ݘ5��"�y�����E�dM�k�|oH`�oȖ��ԦV����)�����&�kÿ����쭢9q���1·��@k���cdrH��h�G�K�8st�=��^�<��z4�(��`߾2a����� ���j��8��o(����˘ab�_d�e��奊Su��Nv��!.�K#�Ӝ�󞞏�J*�H�E[����6g2;���'���"�[�j���(�{#�z^�!�0DȜ�x}����Xk_�(�Uw厕�= �֤�^n����m4n���<�lܘ�W"N�l4����F�XG�i�*=`~a���dTy/�Fj�����<_���T�Ns���Xȇ�}M��v��'=����k>.�5�3#��K��aE���^��7�Hzs��q!l.�lI�,�} D��d�c
aMoBAr�4W'#P��EЀ�r�Ž�ko|�Yj �2O1,?��jC�?����nʱ�}x�� �&�Թ�������uk�O	�Iy`��Y����"(V�1�R�����gޮN�NM��K͛�b�9zY��_�T1���?v:�F���T��$��ӽ�UJk�5��S��R��ӷ�l�%)�L",�ZD�c�GWI[_�l@\;6��Ɩ�(��Ӱ)�oT�Avw=1�Pe[e�lk����S�\M������?�"h�;Ba���ϧR�����e�[(� ���b*���w�v��k�Kic6f"ْ�Hhp.�/Q��E�Գ�fٰW���rr�=��n�i���>7��V@-P�L[)�+��o$��KzB.4�y��Pm����b	�A���]FZ~�	G	*	��O,�)3,T�?�u\��E��b.T��xQ:�Wi�.�W��u�
�t�I����AX.�F#J��{��(D9ܭd��f��aM�m��H���ܠ���?��(i�G�E��ϥ0�&��{�*�L���\V�B��&rajO�X��ܨǖI��ioS%,S�6p����ٝ��XR	!a<:G�C؄H�2J@S�M�O�S��dHEn~��;��������.�@�,���7�x$�cr�e���&���s��~�?��[�E�������F��hw+�	CD������E�vc�H>m�;���(�Ň�\ז�?bι�8�Eͦh��QK[�*&��1��k�/E��!���`���x��"�p�6����FY�N
N�(���DD
��0�Zz;��T97?��V��1�xM�6*Fgj�.=�)O!�.��n�z�ػ��Ta�; ��}z�Z!�MxNQU����޾�\���ׄ�خ�ZuQj����>�S���M]��Qg��!	�S��1:��4J`�d�q���<<Kez����O�4���S�p���5zq?��5	(��U��ak�r�j_���|����;���-��+H±�����@t�$�"�[a��0��}۠�4���9�A�e�y]T����^uW�Ж٩�a�R~DX�q"���+=6C�Ml0��
�"��
�D��%�ZE�pd�g�fR,'��]���'�sm��u-�#?TUF��T�����DȌ5d���w)~�d� ��B�̋���ʉT����[N�%n��S����U��F���0�Ӑ��W1�����IZ9�G���ӄZ1��$���t�J2�n��k��X��H�h)!k<��KR�K���kB� ����Z� �~�e�h�E�z.>w^�h{;�Y�>�E^ڕoTG\�R�H��Ϊ����ɀ��La��*�N��`�Ζ�x;��}����>����%��E>�A���8�J��8���L��d:[\�����n<�Dy���u)|!���̻���5���m#�L�(O���e��:Ci�B���!��#W2*��]u�q�Z*Ԩ������g,������+::vb�t߇�]m���y�7�'}�8%���t����(`�8M���,�57�y�%�6b��"�F�Ӕ��n��g��%�����D�Ʃ��t�R�7-��l=����䃰��G��W��v�馵~�I� �3�$�H�o�,�
�]��J��U%��v����񱦻C�>�GsWz,Y�2��'&<D�:s���<�.Rl�h�uC��l�ˮ�S��Y_�ak��U؟�φ�Y�b!�q
��3}>n�aB�_�W���Z�	?�М�ܿ{Y�P1o	ax�8��m	v�A�[���t������*Pyt�._��� ���v����(%�G5=*�;,�|�2�/Ӕ ���O���s�п���F3�#�z�L��a���'�l��j8��:K^��VT���yS��j��7TA�wXQ�I���p	��s걚�N*�M����/)qZ��oWp���@xo)Ա�����R=#ގ.g��8A���[�',*�[�Tڼ*�
��@%t��=y�l��(b�Ex'Z����K�g���DS
��8l`KZ�8�{ߧ4X岀���-D&�k�6t���)s�694ID�R];2LN�IB�n�q�_:�@_�}�ƖW~\^�5�_�0�A�耑�ֳ�2�|g���we�cqu�6�^O1#�6i#-]!��	��'���OX��x���HG�l��g��|�"��˵� u�~�^��	0D�!�7�W���n��I�nU�H�za_y���F��^��s���=����;%Xhߧ.�X�w�V���D��%V�d����kӗo�bB�k��<��)7zEÒ��^:����q0����.�85$�a���f֔���3I�P�.�>SC�{�Au�!�h:��Ê�t9u��$�Xǖ�U��ƪt���Ss~��l��(M��?:ЈQ�jn���2��N��f�����>> �緝����y�F��S�o?j���{5�dИ���Nw�
,TS?�YG��}���2W����ՎF���v��~J�gK��ʤ�3��@nPި݊���pcOG ��h�i�~ī���pUs�V�%��,�]�`�Ǐ�]Z��Y�9�����:��.�(���[���Fo�?y�ݜ���Y)�����Fl�z!���8�iSR�j����oHl��D*��}��?6�X��������h���j�u�Wvߐ	~C���g>�k�G<�+CS3PͶ���b`Ԁ'��aV���8����<���]�8�L?H�u.�'mS��Y�}�v�ߛ���>���_�cHV��K
���f,u����ZSCv��>f(��csЧ�s�Ag���Z��H� 
ߊcHd��5r���(z��5Ђ;(��f_�S��F��>F�%�t����0-��lZ�?�u_j9�j":wP�}�dJ�1�Pk:6}���*?(��D����D!yn6qf#y��3�`�k�;����ϫ���P�Eq������7����y���!Z{�v�Xp�����- �]71�A�8�t���Mn՝�M�����^i�$��hz(��VM������U��Kuh���򽏎�����q4�x��	�cJL�BG�z ��Vy��]x�o� :��C֏s6�Z��t_�������n���v��o`�@q�ޚb/��q u���`O�MC:��mLf��X�P |݈N/K+���W�2ꀠ�k�O��· `,������k���ۈh��
T���k#pOT��8!'E��G�^?���t����P��/�5���� ��30e�ye�
\ǚ����ۮ�ށho���.��RU��SS
|w~�zxIk'�;��v����B��9U@��y�6��;MPLAzj��*t0c�{�b��0�nyP_Lj�n�ݞ�4:����������" y݂��/SL�(�k��ݯ�������EE7�3��,�#$?7ն7� |�(��xAZRd�R��J�z��h���	�C�k��8�����Q�f������b��
�1j�h+uD�6��i�k��%�J�j��j68r{k
��>��e3()z�<�z�SG��%���χbCmfV��IW�]����C]/��x�v?��klN$['aC>�����^*:z�a�bE�R1��(uB�A�t���_m=�g�'�P�H��E0�x�6o��y]��\���c�AѤu�-��J�+�ݞ3��'�Vh����3�'`��
,����V��?R��3������zZ��5�g<����f1��:0M�tyɡ�r��}%�aFܙ �37%#�+v"(4g%����zvK ���QL���
�m�����4�������o��WAg9�?���^�F?�ɉ[LO$]�3�����{��G���`�BTH�ݪ|ƪL̑4L�z��H#(�Ee6$�֊
����P�J+���w�H���[��`Tr8<:a8I���]i�����@��g�T�6�[-�	���91VK��a�
f_���/��2;��t�Hfh��.ھ�(5m�D�_W�d�37����7z�i�,�H����Q�!�Gw�	bJ��db�J��z?|$�e�:g��s�:��]X�W�6��Tř�qR���on�P��oƠՊ���+h�(<U��o���R`4a��
Q9'䚼Kp��b������L@'���_�s�����5��![��$N�.v
 p.P,�ZǬ��2}":�<�O��(���A%T*pbՁ��\�� `e��;iW��B8@�*�D�!I�	�eO<"D��<z^u�Խ0z�ƷD.G��.�s;��:&v���:�����C��n�;`A����y;P��W2�b:i�c�M�*�!3
HZ��>y4��ʽ$gyc��Ⳓ{��z�f>�
(�j.�eF��HsA����� m
'�'�h�WL���V�7�!�̑0x�)`^�P��cd���	{z����$��qe�8�`��}8�R{��8�}YA��/�5׽ ��|�j�+=߭�����i9֚XQ�yZK�y�a���3�'-����]��ZsOYo��C�)���VC	����$�����vHge�_#�ƕ�2�cq�|1�J'ѨQ�g��-��Я� 3���֣h`%��f4m qkǇ�*k��$�՗w/*���s��� �aR��|ƚfȘܙM ���~'AHO户&�O�R�� �����?M�e������뺠��T����������f�#T	%�J�E�-��8�O��q�VoR&k�5tQNmh[&d3*"͟Sk�c(��l�&k<���E�M�3�����˺&�X�t������n�FLۯ�U	�*��	ް�����U�+K�Z0 ��]��OnP��O8�a�	���Z�@�c��I-fq��<^W���=��W���\�W?t %�]���p	ҷ;S��i,��BA���������#V�'w�6*��ϭ��s_�K�XDk�bE�4�k�l����x�;;��se�6S�5i� �ʯ&s���Q�P����ކ��Y�{̕�%+��I�/fEu�sت�n�/\= ��E[I}��+2O�꾍y�J	�R�����j�mo63D���}̡�@���,�3���hB�d�������� ��JP�[�(�v�w5��K��;��`s�g�-���?y���k�N~��Cn�!7 F�C�V���
���9��;�M�����U�;��c~�Ԝgߓ��9$�����?r@/���DV�z39+�ō�t��.v�c�������9�HX��Q�WhR����ۂ�w�c �l��W��H_��S����p����$���S�,h�q8�%�(�4l oXN�^4�G��M,8Î���=�����5_z��+\�T�fL4pO�xB���R(M��N�->��;�XEu��1��iF�{��fr�?��[ս���6�<ދ8��+�p[`�,�Z��[��K�4fd쾮�p�����:�E��P/�E�4���U����}�z��r��wJ�v�@0�ve��<n�U�&i����J�?'���L��@�n��״g�]w���<a|�W�b��-��!�ǐ&�U��q`z�;�M�קEd��gk�;|�i���Dm�I��}�����XF���KCs¨���;	>���%��댄�W\�I��T��aNGa!�X�ԓr0�|XE�/̎�r��9��/_b+s�� ���+�.��k�J��C�x��|g2w�"��A9l����(0�,=n�\�f���*P�Wh��5 ��.��v�kaP��Z�_�,��N��tR�g���:���1���CT&`���ec咣�D�*��/WO���~d�C�����S���O+�����$����Θ�Ytr���F^��2(CɸS8�Ո=��G���s ��P{�1Yux3���^�o����I�� ���Òвa�[EJ��4?"��RQ������fO�^Ř��Y��������^t��>p�^����C�c���k|n�(�i+��]'"Kr��o�$
dV�а,�_k�L�M�F
���'�3�ݚń�8jϜO�"�������xj�譣�t�K[�̕��pC�o�,����k �`��]wfI�E��-f[�PJ�0�e:�&�-|+�S��:�h7�/|�p�T ��>�B/ypXT�umV�|	�w���= 1�0!j���_C��9{^Ov���Q���:c%0~�Z:͡�s�3k�l�%�U����j��@�'m����^.QO�J++"n 8��&~��K�=+jv��)��6���u�i+�>��a�!m���P"S���!:%Ea���5)$#�|NAE��kd8�'�2�>����6�\T�6y빃�<��|�5�c_�3q��l�2���W�JAtT/�rV�խ��~�h^?�2C{�QZc���Pb���IĬ��z�e�BY��^��f�*6A,����O�dk�R~�*T�Vx,���Ω�u�'+����d[���*-�`��*��N�u���_%��O�c��	ߥ#��˘��U�u�cJ��i��5u��8?<`*�uB<_���iF�x�����Ҟ�8"�t	�~C�iAo��(�(�Q�w���_
����ʑ>�D�ٌ7Άƛ�|ݧ���/B�m,#E��{�'���h`�Q5��JU��M�@��	 �]��f��,wu(�q�{��m�s�+���A!��ţ��ڱ��a<�1����������|�������B:'����� ��TѬ�aCh��X��?g�.D;l�x��,>�h�;������]T.ز9ܖ�q��ɯzK9C�[��+{StJ��1^��4����A8c���Ù<�2G����]���!�<~�{sf�[$4W�mp�G	��|������������X�?�`,��k�a�O7���Q~�Q�r"K�`:5bM?3���[�F������	�t�ǹ��pؒ�㪢�$�9hp�hk3W���������Ɵ_���DQ��Fe�'L�ۯ=�f�:<�"������׻���I���F��EU�S�B���_��J�l�!���P��f� ��hs���g��9���k��6�P�!�G��z��x�:�r�ǵ��2��g�C��Y���Ŝ����	�r�Nh����Ϸ7���-�>�;�CQB�1�YU�Ā��)�mć�n���'V`�[+;��3Q"��x?5���\�x#[���:�d��3B>����5Џ־�5�+ke/������d�3n��	��,�-7�^������ٚ���z�a�>-}s �fyP�ovR\ �A�Cúr �`�u����&���̿1��@�q���Z�}a��UO�����?��Kq/��,�F�q�a ����ܤ_7��z_J��"��!��8P������h�"��u�m2����9��U(�b �9-Mq���Ϊ��!��LVlG�	�� �e��PN�VY��,5���};Y���pRr�M�|�nY��1 �W����\&r��Yͻ��lx�q��:��*7��W�@�K!Z��V�I����E���ְ��\7���N
�S�oc�Ω���+����=W����m>��"5���z� nF9
��[\�}К���$��TZ���8�9�(���婳�,�O���M?�l:��N3`'#�:?����ؽm��搦�,E��eDf�Z�q��a ��#[���0͚������a���d۷I����,�������v�H��Il��ܰ����5�<6�f���K�p��p�F�ϔp��"e9U�i��	��]LVfh�G�	�듧���!ψ_J�+g�������)@v����v?]�P�YVhz��yǔ=�*�R'I3*׭��|>)��so�wv�j
���(��x��b`���l\Q�<(��+>��ߔR/,'s���m�;.�G-"���2L>V����C8��l�~�}�\ �*��Sn鵪��-3*:V������
n�Q~V����|�.��d7���|<B���[ ���:HP&�x�z�>���Ip�*i+^߅19���7Jk��Tl��� ��Beeu��5�)��1�Y �&W�.|��?�T@W#ųB F,�1t+�*E���1�zXWs[�8h��B">C���Ǉ��[ @��Eg��$�'H{1�z*[a�B�+�P�j�`�oa��O[�sb#ㅾa��_�)�	��ȱQ�4�ĉ����Հ�\'�3�D�ј�8H��fJZ?�;�`������Ҳ5 �ӎ9K�J�	�-J4u���'��b���yV��t�o���Y�pM%�\������"a��Ê+�f2�O\����d�������l)�9�-R�1{"'��m?'[)�|B�z�	��<�p0�t\�-8���`e���@�q:9J�MW�
穉Q$��;("�� �!��h��r!GtFi4~'�ˬ�F�d��n����\����EM��r�Qh*�Ǝ�y9)\�����ZE��J~�e/�-���9�XO$�h�yCM�7�*�i��-�-֮��Y��A�=lj��I���7F>���k���kT*H��c��{x};l�~6�B���E,�2s�r��QҸ��i,�t�&�15��1{��]���?�*>�3ޒ�/�.Y��0"�ޘ���̿'"��.�z*�R���n�[P�l�m|A+%�
�@�,�A+�9��@)Ù��׃���%U�P,#@o�%�8�Ӻ�(
R~�P���kK��[��s���bm�&�Ib�2��'�ZU!_�J�`A�����[�ھẸ�К?gk�]�*v�Ӑ���ک��\��m�����!�Jrqp6pe��2&F�0YG9ζ|�c�R�$�(����Y���nzS;6��|VG5�CJO�(��n�K�Yϫe:�� �>?��ǭ�X	��ǽ���оr���;��rIi~
{����AA�k9U����_�pG�rL��>c�0p����Y�������o��)Y�����I�ح�M����;��ћ�-ON� ޴?8��Dv���LfF"�xK]����<����Y3�*\6u�hy �h�����tgD����2�˪�~��R��f:e_����J��.�������]�?�|��Hjժ���g@���btuW���X��|����<M~�SJ����]�8��42S�܅�JY
m�k�Ą����=U��� 2
VU�Dz݆#�����pn����V�Q?����8#��tZ�x�
n��Qa%e����3IJ�
CbׯE�����@x�o�QvUz;��t�S���X�`��؇8�2]�Kv�^V�����O��1�R��0e�H������Of0'DR���^�9Q$[j��g���;����6����F�f��BLF�����`����&��u+e��S�pT�&�=� �>ͧq9�	v(|���OS�Pk�ޝ�M}7Y�0���i�=���-��w���b��CzR�3�ؕ7)���4w��3E�8����m��g[5N�Nl������m9T�3�B��7����ȚIƬ����gc�B��0$����[�ꒊB�#lA��!�/ɃI� ��2��Ud�@oe���}jC�y���&:�dn���Yu���tG�n�y�?��="y������m��n�(���!�ţ����ʚ��[�rwY
2a��_#�ң8=_�97ed�[�rJ�6�e�neR$��'�6�ܰ(�3��?\�u��l贌W��ɘq�1G�
pfg8�F*K-\����4L�Kk��kn��zP�x���99��N�M��~�Y���ل��}+�$��.በ�z���YU��y��iB�r�-<h�52�]�5��jffR�<�k.��j���2�΂��b)��(�g�W��-gL�&M���Dò��y��&H��<t�T~z�:������T���0k�UQέ2��e��/�C؟�g�Ǧ{��9(l/Mr���j"��r}q\�H�[��0�d��2	m}�#��v
���f��Z���R̍�	����k�`Ђ�:"�~��LG��a;k�8riDG!�^��{x�Z�N�wt!o�T؞Y(�*�>�B���t q���ý�	�b���Ȅ��^�?9�_Z#ϱV⫤R�j�#���]�q�.��aĤo��F.���+�&^�̹?�K:���~�m((�j�y9�[����[�`w	��(!^F��w�h=�2'�a 4<��	�5��1��֐|H���Ҧ��`@��䜇��#��'���Uoi=
�m����YJh���3
��n���a�ԧ��]�axS��	
� ,�s� k+�:�+��n=��u�F%����Jϼ}D�ˋ�����d�C�yʂ�p�����x�py���SئLnS[����J��H�W���v��b\��$9 µ����cf�Q�:�k/e$'������K@!����̙�ݾ��%��f�� ��������������KOb�l�u~���,7����������냢`a�\���� D�0|2� @C��g��!)��B�S�=˒˥E�34i,'_3kw���gx���av=	�}cŚx��Z��Ku�������D��q��WX��M���5q:c;�$4�����`F����j���8��w;�S���6������I��L߬Ax=;�?�5��8/���\��K�B����G,���1c'��g\�&U�"ov�=�b����$%�t��B�{ ��x�j�˽A�4��	�1�=��[��C��g�:h����$��4r����=!�Mk�2���s�9
��FS~���Gc��$/�
�V8�vS��b$��8���'<ΰ�M4ʟ�-�0~�2�ԍa��~�K�aC
N�w�D�=��<2r�=��� bCb7��4o���%��fh	P�_YoR\���K�b|���Qd��-�e�a�����<2\��ţy�9u}��'C�l �����Qf��U�;N|��t�o&Pij �VH1eo�ы�7D��ԻS�`��0�j��_pI7�{[��{�yQ�v�Zo�Q��-�������խ}P/m��q��n�5��/��T��qk5ʱ�5�Q��2۾۬U���M{�W[/�������S�Z^�$��Q����^�<��T�ǁ��|?��'�V#p;ǽȋm��`FF�P�Wk�."U�_�x3�!�W�#���ik�*�q�C�n�p�{2�zgW\v��4�ы��4v���B�\��/�V���+�!T)[!�T�_�r�9&��6�0O�P`颰�y3���dV\�װ&�5Ľ]LrN4n�/o���ڷ��S|Wd��H#w8�&��{kć�<n��X('��z�x�wMK�8�_��#�j�9��#�'���4�|?ßk��I��t5�j��R�}p|ö���]ᓲR���������Ҋ%�& �4ٜ��"�p_�ӝ;!n�f�BR��� C測�h��!�X����˝�����c*Y�������|���(1�:���d;����z"�b5܃MXi�]�F.�kCnںCV�R�(�K�?ʷ:�
��o��}�o>�)��JAϒ��Z�S����>�"j�o�B��@���'SX���\q��[��D�6�3������@���
Nq�.D4�z1X|��e��>UK��%&���C��np��%��ceX�����K��⛴0�ͥ"�.2fS�u���F�ƴ: !V~~�`����$XÔec����L�860�;P ����F�ӹv��G�gcx8�J�S��."5?��҂�v������H�����%��VK�*�s�m�v�"-�ul�ہN��C@�u{��D	�b���~pH����8�J�{��ĸ��K���b��
�
[U��ZU�Z��Kz1B�g4��XV���϶ $��8.�Y��64�6�P��n&�U0�����8�)�kD�!�7�$>�X��~�.��D��D]~�1�8�e�L[�@\�f�ն�,V5���5r-dru�Gmj�M��~7m�ϒ}e���t�}#~I�jAD��6���}��W��_\t�P����3��N�Q��� �ɺ�.�R������:Re:�2�H�@�;!_��D�7w���{����͸b���[i���rJ�����q+7N(Ybل<1��G������׫����س%{�s\�>�ʩ��ڗc�X����nڧ�h8��?��.��G�M���ʩ2O�^����
;^GJƞb���8vE��d��Zڄ`��|6�E�/bȰ�i��Y�Y����h��(�Q~�#�����o��wQ��'��ϫ*�ɹ�@c�%b"�q���t��3�O�>Z���
��R�'�ߛ\M���>��÷��	u������׊��.�1���˞�󇐲G�ݞ�Ό�b���,n�ȹ����-^����aX�ab���bA�< Ï�(���꧖v#�A��NJ�TL�`cgc8�UK?�*���m�������ea�i|�r���9Y���YR�+���#N
Efn��,��lZH/^�ťdp}8֋����!�jTc���+�Le3k�EXc6��.�YxY�*!� �i���C�f�`<��]��j^�rv��-����_B��t)�Hl�`��q=Ԩ��g��H������9H�3eQ�h=��QU�z�	
��p�6a9���s A>=`]��I}���6���ΥL!o�Y]]��`�J ��q#�:[nm�EN{������R1o���0��xL!�Uc��h,_G�T��L��_Ⴥ��S���G��jަ�M��g�>~Xi�Y�7��Ug��=��M"�V^�tq�V�!��m'�#p�@�l�zßҕ�z��c8B��. ��b�G{�^�V��&]$��1}�-�l��g�:߽���!_����f����)���\2̍T��1I{�94�)5��M��IR]H�,]�%W�[�E�׌,=[@/HV�j��0�S�׼ѕ`���_(���(��H�-A��	�\���A����"��e��]#u4ʐI��}���$�z K&-�e���D��`MҞ�����Y�b�w��_��������R}�etx�8����"ZQ贿�w0#p�K��\�$�&d�YZgU����žD�b��4��'W�����k|�ͪ����:bB���	���)]	�)a���9 ���qS��ĸD/��G�����5��ZD��|_��˯����r��yRa$:mEi,�b�I���y��;�5NrkA�'��U�H�rG?	�Kp��=������&X=���$�4�$J�ѼJ�r�ԌoZyew��E��IU�5�;�Zgx��)��
���)�y$�n�{���q�%�	���0�Y`A�}M�J ^5��>�̺�c0 ������m4�A{,��#d���+�ِb`o��v�&L���ɋ�X��x��k����5H�v�Q�Z:bQ����EJt�;�5�T6���s�YK���;rp1V?����˧ޢ�?%��R`��ݧ�B�PJ�	n55:2A���c�ܚ"4�f,��r;�1������<�<���&N�Թ>��Vej��Q��]��N���h�m��?�v�v�l}=����Z>y�'4���'��G.]���q��/Ո��A��/��� �υ qXb*4�f G�8Uq2�-e�8��P����%#VȪX
�[���yds��99#�~N��W�:y�=c�	Dtw�l�rc���?fF��EK��du�!���_J4����h	�P�I�욿q�䐛/���YHL���[��tN0�W)�LUؾ��[bV���1~�u�dW �3�������vi�I�3�YE�.�p��?�L86��P��V���@���^�h���� k��� �����2�:�>z���<�/�ZN�p5�
��{���l��S<Z����v	���iG"T��KrP�U2�:�"�g�����X>��A8�B]Yb"�3�A�WIS\��7a���eߖL5V���ί7�0VM���{ᦰ�ŭ�nq^T4c;��� �|��> �n��Ŀ�SN����k�cn|�2"�Tx��`)���y�Β���u�/E�Q��8��-y�ڜ��6��P�1q4&�I���q�Vv	��bD��}�8Hl��l{�Ì���ZI���8�;LtG�|���A�u*P�N��Y:�HU��]���x���i��l��c��>~�UϨ�;�j Z vR�$WN�r3� ���܉���/�ճ��W)
����b⒜����X|��,�R�z=�]�U��p\�i����m��]���� x~��2���DQ�i��e��zW���_TW���Ka0vF�V�!��􃨢�q �A��nM-��P��?&x�ƶ�Ӏ�P��V���W"��t"ۏ��2XQKL^�����-�� �<�Բl�.z>�z��C3]�鰊�lɋ�zb���}l���+��q���Y�[�}=�K����%l7��=H�x6'8$�y��4��8-�T>�8
/l)DS'`�iRoES�����}���WtMW��E]�Ͽ�����Nhb �JKy�"��W�7)K_<�-�n��Y�$�3]z����I�QP&y�>;��цL�(]�U�3����k���2����/�%ql�z�o+ѩ��엷L^{4	�޼GIt�&Ǡ�b��!�.��@����D��#�����pU�B��7F՛8!��i��j���;Z��Y�N�?nj�Q ��[���Ѡ}�����y)1Ҽ��tsMZcT�.%����P��b�+(�\�tOC
���s9$E����}��o/�m�L���X�B�{d?8�əFM�rx�\��߂3�8^�^�ue�D�]�t^)[MFڻ�lm������aEx�%dS�^kRs"#rYcG��C�%͢O���H�bm���>R5z�����Y0�#��2� �r�e,����e�8x��S�^_���U�{^�4}`�}��?xe�7���dHj_���y#�˃Gg�j��.�:�zh��.����|@/LH.'E�P���:��Ndg��/�6�m�!A�e>gWٲ3,7�)Gb�TO���_�yc*�)N9H	����ܰ;��z7w��y9�#���e���Z�>&��0'�CMp���7xЍ=6�<�3S�X�3arh8���e�nE>��@Z�pb��eb�Mノ�I��DZ��r��y �_�9"�e��`~B�)��΁��[�#��8������HBL���RX�	Yj"�w S-�)C�;�7�X���^$D@%W���9y���a�&!���z�	�eCt��J�4mʠ(YU�aH����Ne�Ū�;�u�f�nf���,S>���F��ʆ�rw�~�E`�h����w�C�\��uEI�ʞ�R��W��â���4AWI��
8���������F�a�˪�'\��� gجXqg�Ky�燓W�y�*�UT`w	��E��P�b��M�ª c6��~}֗���_N!����F����C������l�):?��J����t`�� �/r��{\���G�cJ͝=>�FX���0,ny�@���|�����(g�
�(Jys�� )�5�o���y\EI��{+��}O���7�.
G�S�
8�9�U��y����.V����Q(cpd��	ͽ�	�(�|,�`���K{�!�v禡g r>x���о>S=�򟈹C�3��Ɲ�ga�*Z�o%id!�s�T��M5�rUzF0���{��k�th���n��B�	N�3�����.���@���Rz�$���z���Y�O��¦���t�I��^O�9��,"���7.�����K��e~-s�{�Y�Qg��Бd�iBhmb��#��=�2��Jͪ��/���2�aG�|4�`%Pz)l�5���
��������,��n��p�L���ԓ ���������R0�B�B� �R�B1V�8O(�f:�Ѡ���j����5D�0[f��Oh�<����B� &b��=���ҕ:aù%�༉Ɍ�F��n��u.f8>�#r�������),�l�e^��m2��gԫ�i%���|��u�}�:P�A�V��v��c"e�{M�'����I��~�_�y�����v��Qaa�� ����XW�#�<>�\�l~�U7n�wi	�����ԡ���I�|�Nb׋�\p�k T�Ն��,js�)���L��{g��;��'�|=�aեo�[�l�v,��pVĘ#Ho�,�V�=3OL�K�R�P�,��#�zC�vH n����_���"}�`y�)��$ �c��v�@Z�_��v���7r(!q};ưSr��Z�F![}�7���m��lE�6��t�m�6.h�R�aB+��ˬ��݇}H�$��@�җ>��N����癀Is����/S����Q2K�dAxI�~�����yY{�~D��7t�����hS��nCv��4A���(+Q?�������H�a��.���DB���x�;�ֻ���_j�uS\�Ɛ�O���ѳ�Ni�ѣJ�(�y���6_ח)�v#�Q��n�&
�d|*k�>L6u�?��x��Pʐ�����Sj�閶� >}�E���{��7棢�g��4�<�U��� k�0�ac��$��fgDb�S�6m�U�i%�r�
%�Q�Ks-G���+2*�,�?���WtdY�T3K���C#У>��,mn(՗�Sk3�����u	k�ԯD7P���q{���<�M�' ͼt����ǐ��Mh�O�`�Qdޥ�~l%�����S�5iJXy3P����G�Wbx��3��O���8�JV�dy�ҵv�\Q�B�V���]4g����|Q	�G�q���]6$�+��VHl�x����*�Q�>�f� �0����d,��w��!�q�O3F���Mcr�I�V�4���� �	�$��c󒋏�=�/gf�y	��)�\�%P�R��=CtJݙ���#�n��<��ex��po���+%5{�	�M(%�e�"�
�-M:	;5B����n�E��;A�:aiI�k�����G�^8��i^��f5����mD��ڴ5����y>��D�t�d I�&)o�ڵ���h�8�T�ׄB�>����tr����=^]��{`��pK�8s��%^��En��bqRlwB�"��K(u�V�M~�:ҧɅ�_̈́Li�签{>�{�����,�w��S҃c����<���/.�4`� �&�{���4�y����e���O[/NF�8��c����f�G��&p���1���Y<��Xb:��K#�c�:�dԸ%'����c^Nq/�_����lw�/��^*�k���r���%:Ꮄ�1��t���L�{A�(�c"��S7j�ί'���.���U0�ś�B`\�Iv��xEA�)U>{<���� �9ٟn��L*`"^i�N��9T6���kn7�wz(@F%�9?;�Oc�9�i��E��̷�S��ꯣ^���Y��y9F�����>`Y��E0�S'�*h&�w��*�O�+֑į����R�}�Zs`X�m�#���g뫍����r�?K�b?�9��K�1���ʼ����󠃈��=�z��9S����Q�YE�O�0-��"��a���;d �w㜱e�=A�K��WS����攷2�B��,"�d=u��RB��"���>{NJ��1̶��?۷NeRծ���2����Wh��rOM����X�FP��ur��!�:�H,2�X�Ese��0՚BQc[���6���'�$�
|G3�����QŊ��.lv\��FS����9��=`�]����~�rz�F#���3����B�Zt�"��kৠ#�k}����djp�����P��a�4����5�w` ��j(7$��Q�ڠTz/ �v��Ai����K�?��l����*�P���A+���68\�Z��V�[#Q6^y%B�������p��WD�N��wׇEN�:�+v�O�"ۯgx�{>�@�(��YEG�.�4�=������>�޽3�q>Bj�<�g"9�-����/.�-�s:�w�I���
g5q?�U��L�+nj��(����C�ܤ]'tBި���`�fW�s%���R������ĵQ��{����H�Q3%H�z���O@��yf�Mx?�ďo��z,L�S�(%� \�x�'	*Ͻ���kd��QO�!D��B(l��2�A�2�T0[��S�+b��=���'>�['���U�Osfy9H�9��}#�6	�IU��	s���)����>)� ��}1l�V���<������b��'c>�����W��q�I���q���3u��I]�4b�V���rEć���fF�tηP�Ɏ��M��[��el,�!0�t:��B�6�`�N1��6d���:��Y��o&4�7p�_��$+d�C`U��|P��b�Wm��P�����̦��zn�Ov�C8�kM�4�G!�Y��_
[`B��C8s
��[���EE��vz�$������'EÇ��uM��E�,9�Z�9��w�'��~(!Fǫ���)���X����g�M|v��J�2q�h�bO$��+>>]��$�F`�_��{{�S~��L��?��7�C%���VL�ۗ���9�^�m;�.&v]�|m� 5p�s�w�n+#rmE^7u���f}ϴ�&��CP��)��@���
�l��U�|�B^U�Q��o�pP���ff���6���4��@�~m�f����x�rz@H� ���Y���a�Fp�( ����d���w�Ċ��!�y�Dc�W��Pv]����F�h)qVd�W�VZk+A��?R�?�%ȵ=a�mi�BD|��"*pIOP�~��=pB�q��J�+����a�f~6d��&�)'k�|9ᢒt���]��n�H�ւ�0��-k����R �?7t�Ϟ\v��b$�=��5�N%��zY�����#gB��2��o���T=Z��4%��#e���7Gl2~BZ���!�Xb�i]VM8ΌsQ�%��ICM��&i(T\��b��S���?6��}\��*%�ܬ�֔�`�	��|6��P�J:V%����wM~�Ȋ���(ܤܴؿ��z/�N@����_����߅P�y���-_;ۊ��b�o)��_�W6���cL7���m��]��dD��4:Z�$|���z
ד��N�������\�,�U:Pv�����mZ�,"���+n�r�s�|��]~�6�r���U,7!ʌ�}z��_p>��*Q�#�<��̭��u
�Dxk�#�x�;�8R$�w'	����D�j�1���x���l�_%KvU����W=7��U���te��{���V�������;{�3/��& ������ �A�U�M��$��Q^��&[����o�n�*�C������do8�9�����/p\7���t !۞���䗢�࿐:{�����a4J��A5��Ӈ)Z��\-�.j�nd)����nK�So�'�&�t!�)�O�
E��W�eOHp�$ke9��4�����"K��}Z���ʉ����"�W��]�_�H� Q>3$�a�?5a�@{�+�m�3�t�d�� '�y�~��/�5��q�n�/��o��6K� 8�_hM>g�F��c����`H��OA�D���h���>M�9E�t4rZ���gSS9#zF��@���%��S����"@��TB��JБMVie�$g����n�gΪ�t�?L�����5�H��ɍ��5���c�nZ���L���g�Q	��,>��Y�o�T.�%�jH�I���
t���������7̌vw��J�ќQSUҙhQ����:n]�ς�X���?�0}��e����w���\��uW�U�����R�*�]�bZ	����XmPϘ���	�HD�2V�Z��X�\��\F�Ȁ�~s�kAtq�6ˇ���fW�0��x������v�%�g���ʮbX���=�i�<4u�w�o#��lE X!��<#1�hoüxK�.k�\�����!�� �a~r��Nm�T���2�.��6|ߞ����
ý*-���[1���a'2t�Z{���o������a����t�=�#��$G�^!��������YU���gz��i�.�n��w�тg?S�&��m��~s�0�B��+��i/���Juw�� ��uD*�$)��젩ʧ4Ѷ{�3��i�0/U�~Z����{N�|�n<���C(GS��@�C�ua�ǾG�TKb�[�I"��� .��i�;頲�V��T������E@��*�39f�:�w'�/cE����&�.�`L�������1x2N��&�J�b����r��"(��Jڼ-rz����X�v9 Ƀh�y��m6?�l�� �Q�b�������0��DA%zi��s����=Ω?$%o�lo�06��?����=�BCteC�H�1a���wV�ė�P�uj�6i}AxPC�Q�C����lV������c�V2=#E�����Uё�23�oÂA��9��haJoBe�J}���{E��~��G��@� o�F���K$�X��IM�#��0��<*i@K��b����5T��t�C����Q���&�Z��{�f���q���� 'I	7�u��-�����_}؏dԤP.쀠�Q����f-팭�p��tyx�B��Ne�y=�I��1o6& &�V><����/B�E)�`����~--~D�U�ssy{�ea�R,PJ�d9���-V
��Ə�=>�v�F�s5`���qp9��{�K�sL^VZl��IP����h5i��%���5
�p��J�5�2F��N$��Hא�$'��<+�gc��e��?o�[�{؋�q�9i,B��҄��ёo�]���:�%1)��ڇ a�Hw��h��;�f0��l����-lc�4M�=:�_���r_�X��즚ªF8ީ�9Jr"��
����3I��X�.��e lY�,�A,��`>�2�Ž�#X�r����Ah�	 �6�vc���EAX0ޢ:� u�"�	Dl-'�Z~A���'C�����D�A�p����~��k�G�Zz�@��w�OW��,�ʞ]�nͷ��C���Lo�J}�+fB�?�K�jj�R�E��{�(:Lc�A��ę�`W���fe䙆�w�x!e�m���'��~]{udM�lIH&~7Q�r�<�d���(�>E�F�6�P!ȇ��~�R��v^7a���*�6�.�ca*����2^fq���Id?�:�_�ޙ�A��7�0��7C��;Ʃ��3��j7�dx�f�H\Q�|���ɦ����D<��y�� ��#r�-1�l�+�	5���%VSx��$�M}S�Je��:%���s<c;%�}�	��S�=D]x8%!�Jי:�J��80�N��+�i��z���	z���.�-���o�<��=��G��aGf��{E{�Ҵ�����,j {F͆@�Q���o7���BS�� �Hgxb-����TE�cm\gO��7�j��qĘMs�s���s0G�B:�� O�4(�ڔ���׭�p���q�
c�k�Sp��rW&e@��N��}\��+����Da�"��-�"��\ʅi�`R#���T°������#=/���]ň�o���d���0�Uj�$?���f�r~�����,��n�@�V�oabѤ�@� yT����"����� d�58}��dck�q{���I[O�?k)1U�j�A��`�_#O�M�E*�V�!g�8�����&�Q`!�k�.{̓y���T"E�+�Č����P]>m�Va{ .:� l���S�pX����t������>�aU1o�R����~>Yw2��5��@�$A�>4� ?�� �4@e�����Z	�)����A ���RWR0s��p����G����>��p4�BN7t�{]$�0��Q(]A拉�^	홦<Nfx9����ə�Ь�]&���%7��J������q�1��(�K���1�m��r��eܻ���t�R녞�C�鱭��3��Ҕ�&}��Y�;/�-�NA��j��ލI�i�4��E�����լq���L�ʎ�es�����+=\��0�m�݂��,�?�ϮP�)h�1�Ѿk�끣��,|�k������H��	�M�G]	����.Sx�{Qv�s��xے�K P�&��P�%Lc��a�@��h�s�`�v��W��*>���Kn�C3�$L���(b)I���sP�7��T!88\��6(x���Ƴ��&��V�6I�t��w5>��5�W�^���A��_���װUR���"=v01�1&_z�����vͲa��0[Έ�.mѫ7��e�9Y�RyX�ؾ+���f�/)=�VWm9潲����.�͍��;��\��/)��nR����,�1�|��}>�����.����q6V��>ۯCg8�"&�_ }���:Z�,�u&L�	�˅?9�R"���MN�����rez�ԛhjEx�y�ff�$�_�^�;�L͊{���\���U2yX����d�ݖF�C����=u�:��Q�6'1���lZ�ܦk痒O����n��Dd!�3 ����F��L��M]���4�� �=E1Ղ�bgh6��q���I�+3)E�����X�2K"�`���i��Rqq�8���5"��O$$�, �xZ���Z�<WKZ3�5�4��{�~�G!$ ���\Q���EF)6�,cb��V��}F?<�HPd�/�W^�q�$6b��?aa�MN��u�g</hz]��� ���/�՟���B�d���7;�<ٮE� U8�K���������<��|Fs+������*/�o��1E���,�t�W|pp�A�,)p��r���3�#j�z~�"�ȩ�r�@�s�U��[;驗�Y��EP�Fg`N\��fx��y1�����CT��VG��)���B}�K|��2��f\�9�����h���x��������vZ�Q�ͣ��z���/�h�і�(�Py�֪������vYqy>��\�9Y�|k����/H�F����c��8$hK����R�މ����=O P��o�L��)����v��|���q��WA��j���*��&��|~�����צ3J��B]��'n�Q6 ��I+.l��^"%�k3ErA� 0:�F��8�J�ΰ=�6LFld;;��귫��?#��C���m�-���/��ő�d�� (}�M���;ɦU ��!b�T�UI:�l�.�N"�<�Ns�ߡw ����FH�Z���;T�vչW�L
�ל��S2R���aL1����L���ˌ[��r>E�F�|�@"�LUU.�k���1t]��*J��/;y[C�Ǆh�ET�C��fy ���gy�����6k>�UA�"	)'5
z�Pg��^&#�fH(=��/�f��5<�D�Q�_�TP�H8~���;c�ٙ����3I5����D���
2�'R��Y�t�nX�cIq��Y�[�9��b����%G6R�t�����,��dw�\�a�f��^���a�k1�t���/���a:S�@��;���H���-��m�"ZN���ʺ�q���~����n?�%�Ù��Hx%_׮_H��{Mg�����|/���:���o�"���*{��h3� �ܢ��+bn�dD�?��T�Z�M�}��91�����0T�Z<�p�:����m.=qρQ�<�Q�uHH[�D���^�/,l�r� X=((�`��N��:s���Τ��~AU1�K��	/R��}�w��AKd�!��c�+�w���|�߽�,�����������~�N�]2ُf�ޗ�=Z?��ޓ�2��jc�:n:�rq-Q��������$���} ��	6kF�!���������C�'�e�W�>yS�0m��Ʋ�j��؄�4�#)	Ի�Yq�
)#��JS1��R�1]\%kqDS��w�޻�V�cSMW(�q�1x�sG'ۧp��|K�<�\��`��lԊ����f��[y�WS{&=S�
��a/"�!���,�CW;��������wݳp��-���NwOP���
�Z%�^�#ɬ����T0��=l7U�0�8�#)�����Z�N�/� 7�u��dx
���[kV{wi?q��$~.��:?-sPK�&/B ď��bK*È`N�6��	a�d��~�-�t�B/��]�m3���'k`���у熡�N����Fq��p�w6��i�*���K4��C�bo���+���7E����Yaފ��{3څ�ayc"��be[�cR�gM�_��ng�����U��B�?�ѳj>a�&O��f�6�E�^�_E�����v� �i�F�����L�	sp2���! ��6��^�,-���t? ��Q������P�Y1ƓYg�hK4�����WP�(X�J_EQ�`��f C�X�ȀN�Fo�G���N�������.+���u9Fׯ�8��bn�P��TB����ۡ�-��KT8������y�G��=Q��sw�t�њw�W6��v%%]�z��Ky��ʼY�p85\h%���Z��-2�����2�5N�Y����$�+�=����M(�r
�&�v����@�\��i�io����>~�{t�zK��5 ����F��n�O�gM�>)-�5��������,��}�<5��tR�a9�탱1rQ��E8y����s�~ ʳ��,Ϋ���.&��*�wK�Sü!�(j{�3Qlք'���#hoo�wZp��>w�w�aE$R�@�"ƆW��|F�JL��
���6	P����SP_b]x��x:��В7��E�W� ��!0n�~h#`����Ħ�������rJ�@�Ao.�Ν�b����/U�C���U`B���L2i�٥e��ŝ�T�1E��3˽$|�p��S�U���@KD��t��+a��AD�6��j�:�`�3Rh[-�$��4f�=pv�	�e�A�j�����׭��BhBD,���`7��� �3-�b����4��,z/٪�8�7ģ��˹���^ ~���x�v���H�{�Oz��Cͳ:��"�Ώ}�_�Gm�D�,��g'+�X.���pu��uܞ�YCmf�[���rz����6?�v�6\~�\�Z��Q��@_4ub�b|�e������q�2�H�uL�9-C�������1ţh k���X݀�Vǫ����8�&'��_Ow��ѝ�9��zv���P�˿�Y��VKaS�Wc�)F(����D��2�lS�I����"7lJ�	
���g�����>j
�ח��F��]��R)��=
�;n8@c�"�_d�����Һ~�q�t�$�p=�S�-5([�l�эԂ�#h�6܂�{"JZyP�u���YX�<�~}�bl��܁s��2�u�Lnz7��|���iYS���u�A8q$Y��j����6�/y�Q� \w�m�K!y^(�t�1���POj��[X�w�a��]�,/�?M�����1W+��ӛ����j+7)�Av� J�w74��w���:;*L��K�r��I�H��2������3g����bR����~�u����*b�l����}mQ��0k\+�@}�U>����&��(��5tC�3�j�7=3�L���7-+c�s��K�}A/6F|��ܜּ@$'9+����n_y_k��k< �$��^)e�$c�N MG�	��
�0�X��~��B�~R���ñx�Y?�>P���A'��V��sz:��u$u�<����t1�5__z��eT�	�HQ%�RO1a�q��`�<��n7l�7�%: �[��6��"���DNg�2͈��!��&�^�=:9!1]:��	�Ӊ}��o��=n��Y\jeFܐPM�fKa��yC��ڵ�L�ee�g�O��/�3��h��>f]�W����N��"���Сm���]=Eְ�7f�(��55����PU��
.���ʶ��i�}�~r��� ~=;5"C��&���+&� ߓQ�7����[N��>���R�n��ȗ\��о���qĊP�&��P���g�P�Փ�_<�Ϙ�/�{ݹ��Xau�]N1��=��v��t8�eO�ѿx�g|#,,�pӡٴu�.���,6P�؁��q5Ї@yG|<�k˸�H��@)W��<d_@�*ݮa���۠��"�	�aɋ�Ć��� �G𣎺�ʖ�9��r
�O|��A��B$%3�t�1��d(j���>S[�70R_�}�Y<�	^�.@���r!��}(��Zw�N	�n����w��7u�=N[R��X�'ǳ��K}\��JW�����v?y~(���v'{�
�WI+��Ë�i��;΅�
 ���dv��ߦ����Q\W�B��&�+�T�%v}m��3E��1���ֿ��j�!hT�"����/:��P#b/�ת�������:�W:�s�G��������(�\�RLr(g
���'�pm�h�w�Q�� �u���������p���6M^Ա�1cds3�s͛��5�QZnUL\	}�k���l�#u#)E�P������ö��E�����<�M._)�ofs�Q8:�U3�E�
�`jT����A�H�<�y�G㦿:pPvĊ�X6���g5\&Nā`�aC��׹➜#�'%�g�'c�Ŀ_s�x�	����^�5z�Q��;��(�o��ʛ��˪��7#�yXx��5�z���il���+����T�P���3<I���F�V�iA��T��*�
̶y ��K\���#��r����Fk��G�EY?Nθ�5E㷖r���Z��?��*������y�%��#F��/v�������^m�7iѩcҹHp����`����_�m�coZ_bzn�~E�@��Rj�5wy0��E*���Vo��E����S�ۤ�����PI˰�[�Ւ9���@��3I��T=�_!Ӯ@�!~'�qF�L�V�"����2���¼���$���;ds�ӄ#���;���k�{�d;���|9�l��p�,Ģ�B*uY�Ϧe�JF��7�� PI)o����7]$]��W�����^m��oJ��ΰ��g�s�KX�Xn4|�5��~O��Uu�#�߾,w
r��8�ZUR�C���\-���a����*�!]���O���Q�\V54���Ea��0Sxkɣt!�q�Q���a�rТV��S���@r��l&H�p��ˌ�{	�e�LH�����f�q3:��3:�ښ
���)I��Ϝ���� B�7Ԇj?��ƀޓ�-��ʸN�����7|���� ~�9�?w\���������̽u��ɷ8���C���>�3�3m9f�.�jZ��`���<��	�J��*������	+#N�Yu��\�7S�I`}���ȒOa�
�%�V݅u���	�o���^����\gѰ	ܾ�J�09S녶�J�*ʩW4�m�F���6�l ��<pu|1ga�!�R�;��c�����Af�gX}�{��0�Qr��s�:Zz5�eD��]�.���a��!��ѕ`�Ww��)R\.�!<y?�о$�8�ٔ����N���7���肍��̠���2�7Q���0����ŀ^>�[Q���h��o?u!Wh󵰾T�\s�m�&����}b�S���]�ntg�%Qx_u���X}��{�O�ضi�f����#+�����|�ٷW�kH�5k槇B*���c����]�(��N�U�8&�L�7������3����sl&�L�`���/*�
�>�12��d���U����ԏݩ���VNq3��u�=�8����������Fxv���+����|V9-�dyJeHf��1�Ӓ�.:��9S-���;�YR����v����r��;>4+-�LF��<�uwD�9�)~Tx�+H����\[�v�Kiк��7��Ҙ�;��� ^���1�SC��pm6(�DD�%),���^݋}~��4�z�u�~�3�w�h��K"�_�A
e��>P����wC��[��?�%ye��g�Hv�Y>:�j�8�?���,�e��$֟驘 9�����B��ٛ"طꅌC�s��@�J+�m�+�=+��.W61�da��c���� &V��Gotm����� ��z��;�Y�­����{�pY��~��S��٭O�����/s}	�Z��p�W�-�Fv\ǝ�"Z��h ��F&��E�K��VBa��ꕿy����M�R���v֕ꝺ)ƛN-״K��o���*�d�Z��k��Lߩ]"�m�i"���L?UO�����l;W���G�6`�&�=�^qE���+��D���A�+(C���*��7��3�Ϡ1Z�p�wgԂ�Ґ�yt~��(n�U$U��f��i��k�"��Pz@
�=O�Z��<�d��\?󀓫�s?�hM&����w_�����W�x<��ӓ�B��Fx�؂:5I��;$���ei�t�=��,��G�7�L�:���o�;��2,&�荙4o�&�f�i�F�m�e��ɲ�m#��y��yx�_ɀT��L�TD��;!����D�	ȾH�a�~��鳰����rIဟ~*�I��k�k��#>�_��m)��-^n~܋������&+bd@5�d�n���VopL��g��>�ŕx���Ы��ڏB�;
ƭj����]�t !6;i)<[x���F���h�q�O��n��Y�K�#�ﮗ�r%��g�0A��	�x�@ bNwj�����s������0�&3e���&�W��;{����!$�u�f�7%1T<+�����1����i3��
S���L��Ͼ�ٞs6R3�dW�<l�D�e�o-��j�Q��Xi;��xCP�
�(>�j�@�y��C��N�xm�Č����w=�!�=#t��,q�wh�LZ���'
YqAC��(*V��3�#�UB��aO���Y���B�E^[qz�sy�rJf*��cg�!ݍEtP���
�b�>0q9�Q��K ��)@��T-K��Nk���fڔ�GVx4>�\u�K�-斸G3@��k�ZL��,�>g�%j	-6��볖j\3�}�0��$ui�N�k�y"����h��'S<�=�<���FBXi���I�2A�	����`���*S�;v�񆂠�2���b���+)��0"�Z��,��kU�qF���?�k(�G�� ��p��/zߜ��X��"�>0f�Z�F2U����˃X��΍*/'�j~��@T:��>��. X�g��M\��}]����!�5�1}^�,�3�4G�f�#�5� �)yK���b���lo�����R��� ���$�U�����|iBɄ���2��u6��K���Mإ�d��)K@��EՎ��K�?y�����G��檁�M�jl�w ��u-��Pz'��;��I�h�(tV2B�ҶmV'���i�uV����z�%�-�D�L���D=��u(�2w���p�s��?�+��M�u�A:W
n� -�T�@KU���"bI�J^�T�zQ���r1~�w;�2���c�h������Ny�	�\�:]�]��u�+���7*]�н\ �ϵi|���*�ьJ.��F��R�<8�9Uٚ�ޡ��PMOqD�#�F��[�B�,���"�ҺP�K�&�
5f~�F�NO�wܮ;|x��J��k���lB����+�U�A��{ݴ�C:��b�hC��ъޏ�MƽN���Q�/�������n���| .��������o�M �5���D!z�A��l��G���,@V����>;�!Xu�*W�E� �O2��%��Yc]0B��9���~K=_FA^�_�䆏�Ch��F�w�o8�:��	Շ׌����U����\+bY���UjW�$��n!��![�A��˅͑��D��Jq�*O�ef[e3�.� �`E[�,�g&��.���py���h<��6ey�\�K��i,)G۔���ȧ���rR߹,ks�$_�`�1UϜ��Q҅i�ǟ���[���������`$���+���]�sq]�{;I�d�I?ʹ��GX��3\hiegFp��mUS�U>���r�=���C��:�ʼ�b�b3Ҟ�$s�,��e�r1��x����kN�\���nX��u�������*�9dD�f�bl%����%w܁�^�$B��.j��Q̰׎�����W0���]t���+��'�M���U�bΨ$O�5T��A<i�����cIj�{y��� �<�B~%BW87o���r㼢 Mz�}�V@��!����pͤ�4�7u��]�,#����Z��0g3w����qyNpX0�u��[������xn'*�BD櫹q�,k�R]4M��&E�o�����Jb�ޏy�^�]���A2*���g�T��ϥ��(�m��һHˢ����:'���tw)�� c�����4��>�n: ����9�>IPlj�;B=�b���U���Ƥm���D��>�瀬w���v�9]�d,�#wz�a�<À9w�nᆹC��,���Ȓ�j�3�ßH>.�ZY�+o�7e¸�/�GZx.�b��>��)�����Ts�6�&��:�l�,Ѥ� �K���+��.�z�k�S;�l�J�r�W�ݵ�ڢ9�?�/�[7Pun�÷r�l�.�1u�9e!���=�*E��t��r�~�-F��%R��V�6p���d5�뽌�4D�{��^�AD�N����{�)�����Y�y­������biӖaIR������fU�����ӭ�@-��L�_(��T��|9�!i��v�(�>���c/�����Q33�� �T|�;>�6�G���" m��2D��	k���;��tJfm ӡ��;
�mJ�fa>j�� �9I ��mIg����P!���i���"�NC��@ز���ʯ��3ߠ��;b��$��tԂ.�0CY��l������f�뚿�[����qUƵ�o�*L�U���)G*�F��*���Q����V`<��TO@���+ݒ������)vԢ\P�"����@-OF�&;��It�7�\o�;�t� l���H/�.[xx@ɚ��^8ܰXN�~?��s}��F��ʎc�I� �j���w�m���)�-r̊�����}��!�1p���g�00 :�;"��A����Z�p���hu��� oB��D�Pp���A�Cy���1� ��/�~�~ag@c����)fg���M�Q���䦳y�i�̕p��z��E���3�26>|�-,��� GI��j��_���]�`j�m�
';�������w����Yo�XAgI}���)�F9���4�)��3�rY�:i�g}�ՑH�E=y.���A:e @��u
;�IN�I����"t��Gư�sF��N�t����9�׵��<����;��}Ty���d
k�~��x�3�ȅ�ؓ�r�'% �m	e<�vS�]�R*0�*�(�o����V%?�ĉ#�ۚآ�5L��ZKT��*�1�˓�s����R����� �f��L��)Sg֟E�ϝ��Ah���c��㫗J��G����AV��oud����9��Z�J���k��� (u�Y��'M+�2j��i�����+�1c��Иk����.ܧ�-(�;ȗa)hSV݂{�ޫۃ(RΠ���e$���L/�S�1���1{�L���x�m�i^�h9ѧzV��˽ �$�(<��mKy�7��&�t7ک�����A`�^P��kϳ D��]��D�O���#U���@��5'|ɒ{>�r�<%#)k�����<�����hf�%��BQ������ָ�4�b:W���<S�������.�FC;,��H�%~T���}8�8��Q���ߖ��� |Ჺ�"I�5�Fp3u�������+�KQ[A��^�Gw)��8�m�N9�~_%I�Q�?¬tN:���4f�� P��/j�~Ķ�^B��X��5V�#eCT`]�(	���m���R^?�G㓛�YET��D�4�Su�v�S6*�m�,�,�����v�M��J9jl��dr.�h?,/�}:|���B�B�K~��$��dE9隸&� �b���z$��S)����5w���){2I��2��
�d-���p6ه�u��b��*����fA8��<N(�}���6.�@�x��gPYHr#ͱG{�Wa��i�_T�S��߆��@��t�Pm�U /(p�4h���Y�J�*��l
���kq�Dǀ��i����vLA����L�;>���9I�;hk-��
�Ӛ���ލ�b���B�*�%�c���_%Bɤ�5�ؒF�<�B��';�:Բ���ܼ90�x�%����-���E�o��'aZz�������t(�D�`NG\}�j��u�%���ť&��4~T��y)L�� ���s=�)j��nߊ�]ST��ʛ��ޕ� 
���<�y��dd*~v���3�<�T�ƥ�-d�qSh��t��odC��\�y�'b��o��Gm���1�.����䩽*s�v_�5���@�r9�}5 ���l����O������UgD�D�$���$
�38���G� ��4Rb��V��+�b<n��������|zy��Y�����0��	��A?��|����j���@�bw��T����>߬� �S�0�d��y�ʤ^��P��e#�n��O���,�JK�Cc�	(�����^h���6]������ۥ��\ȧ5��H��&b�t�{�� xj��?.�|�������Zg���������E=�|F�	�p\��%/�4��7Z��e��:C>(�vM�՞��NlP�^��exr�!#�_d{']}k��<�v��M��V��a�l�>r�.BE�{���/��3����K�()B��h-9��s���{�+�9�*E��5�tV�7�������Ŧ#Maʝ���R7�W|I^�+����_��J���ͪ��nkkW/E!$����$uX@�#\�/Y4���eQ�;��#��e���B?��D�ι�n%�N��nXP3eE�.�Sã]<�\���HCw�%��5US%��J�xؠpb-`�± r:�F�/��C�N��l	�ٝ���k��9���R��v�~y�K�@4��K*���g�{���v��z���\�j�H���P���$3������+�釶N+��8��K�/D�r!����z�ԧ�Č�k�����XӀ�`=P5����!6XS��3�C�$G1���$F���v�#�!�B�H�<'Ӡm��������ⰹV�2S0?"�әqQ.���I���n|2���� �iq�����$4�!�$� k	d6o��U��^�l�B�y�G�Yd����&��\�= !۷���Pr����;�l(֜���t��'y�h@y!��;Kū�7�
ǳ�ܴ�[���?�eU�6'l/�6�I�[w^�jm�q���E<��X-Ǽ�j}�)Q��5>�璩o���!�� H��GL�Әt�zx���2:��$6Id�������`�K�d��RׂP���
?/��k_0#_�5 ���
������v�T|�]�ǹ�O"�.:n�RKnܓ�B7L~��˱������:�~�Q�c5/AD�
�܇u��va�����\��B�|K��n����F,!cY���h4�zG�Z|�����s$��(�����w�4+��������49H��嶜���1�r[�vF*��e�F���=#4�f���aT��J���֞�j`ߏ_Nݒ	�U-P^E���3 	����
ps1R���I���|R�\���U��L.����h�a:�f�b��ُ�ك��̹��[�8�%rn�r�[���y��p�GS9�шܒ�^�pj�є��:hC���y%���RAi1�["�E|5�đ#a4o)
A�Ч˫!�p�%�A°/_���Ռ�8��jڢ]�74��e���÷�eɗ�	��#�瞾����	�)=�'{.KԔF�����m߄�:���,p�|��OV� 
X��J���iC��Ȫ��}�6u�J���D8��kC�)���(���+L��*K���T�Uo��m��K����=Q�DJX��U��)d+������l�yZX�=9l���½G����L#��Q$,���� �A�O�&���!L�B�#�Akmّ���5��O9��7P�����V�{Ahw�&u��P�N�O�S�BX��������y��W�@��� 䋞�f4��7�a�����J;8N�]��X�e;07�lhq�/��5�М��H_������R�x��W�lL���ޫ�p����뢷��a>Ar4��)�HS0��G7���e�ky���H,�CQ�?ۧ�IF�ER�z�ia�⠒�a�z�*X�]A7�+�	�,����b��v1P�y�̷>��0�z�.u��ܲ������<�@�5.l
��,{����.�/�Q��z&S	"�w�kX�FD4�P'��|����I�ii�3�ֳ���c��Z8 /.u���>�4��R��C9
�;����}��n\:WD\�+v-m%i�/�{",��%)0���oR�'-g���i�0��=ky������G
�FOL�Epe s~��}��K�}�.*��l�aْ�����#��n6؟?��rBq��?���`\�K�ž����[N�+p�q����'��0[��I��(-�#`�q�1X���c��,\f=�2��%
4����ў�g��˓b2�
f��'\S`�/[�[��)�o5d�#+�HÃx߁_n���o5 ��b�0(\�'ʐ�>sQ�}2vݷȹfl[�1H���"�X�Wh��&5��Z5�DE��$��٘4H	g�
<Z�7û���5N�M�@�- ���ڳ�$�VkPc0�k�_OeL�������=�:m�\���P�X!��=���>�L�0d���S��5��2��QY9�w�S���Dm�h�W���1�7#��wE,6cx��s&��s\��Y�����ۓ>wH.2�T)\tz�E�3��'��C��ޏpz]�O����lHȠ�'FS�؉��\����ݙѳ�-J�����+"��S(9��������޻�zچ��UU�-6!�CW�ll�%mN�\�^!��32d�M�S'e��փ���2���@!��$0>�������YsFՐ&1�_����H�N%Aֆ��bq���z��V� �|�2�E}��hnMp��*0
)���f�]R|� ��֠�a�l�bz�!�zģ��ڀ�r�D3|�6'�2���Bmנl_�6�����y�֘��	��0�v����9=�f�an�kc�~{�x�\{�[j���,��Z��8&��f����CN�1��-��V�,��Ba$
�s�H|��h�<�0����q��Z���J������ E4�yk6��4[����zzj��{��8%�2b���^>�`����n.��K��u�ܪ������}@���B��@Ƨ���y�'~��Z�*�^i�Y��Nzxګ�@���������*�����V�uQ��QF��Sm�)����$����	��姂�vh������'Dp�:H�Uq� ϳ�}l��:��Y:������*�D�F��J�\��J3�ؤ����4���0���T	�e-=���0�Q��Tf���s�iоI{�gZ�ݱd`l�V�Nh� ����m!}��→D�Q�}��E�@!��]1u�&"�����YA�<S&b�w5dK���yn�\2f��2?}zUwg�Vf�6����&S��J�D�O�3�B&��0��i�U[ft�KTR7�c:�� x�RUr0C|�g�NoR� ��Bt�M|A{KP��/=)44^���������zK�H���i�Z�bHy׏�����b;;-�o�0a��B�JLʾ���mէ���S����~]P����Ȉhȭ哧��텊~�e�qE�}}vm�G���P|�ߙ�\���/[��)<�͡�mN�Z8/
�{�CU埧/���X#�K�8M]��0���ӊr^���/=��Mx��
L Eu�T�ea�r�j�R�H��)mST�4�U�J���!�F|��3�-����,�[���E��6:~��b2��:ը�^?|m�&ۨ �E��^�
�Y6a.��Ɋ�mH��ts+��U]R�`㓖��j�P1�6:�.���C �V��O��~+� �L��a����4�g����ƺ]��c�Wr��y޾��V�x<?���-oј� �|�w�s��gxDS4�w�Q�7�Po���$�f��IID��	)���v��A=��
���2��3�����u}��2t�$��}Q���9g�J�Ao���U!ij��D�S�����?}K�O�¦`��'p4NU0����G�g4���<�+X���E�
D�_�Ѩ���24�����է��(r����T]��\�_Jb�3r�A�8�Õ�_"�!�ax���-õ���/	��k~�t��2�� )�nQZu�ի�H���P>��U��hr|�!�o���0�Nf�63pp��7�tm�'��5j�����e�O��p��P��o%y�h��%?�ٖ޽��0�.%��k�<�	{D�a*[��ߐ��m�W*y)��h��"��{$DN��3�`~�ne�MMQ�AS��Ih��V�?]��Mu/�Qe�b���k�gQvX�bu����("DO1C�	����-9"��(�T�c1�B�vr¯f�΢��e����r��װz�ҭ4_�������ʞlDp���[�&�܋W�¬O�p�����J|�Nj�g,\t4V�)RVsY��A%Q��l;g!"�F��`1.��i�-Q%ʑcd\�}�H�xvL���|9p&6�Ubl�/�.�+�{㠭S\X��S��GE�����ҞUM�����f��=�Lb#���
��U�<��O����4�c�K�#���j��b/84��Վ�:e�Q�D�ߨx�E��Dq9���f���x;�6З��@
����X����4bl�C,�K 8C���RDZ��&Ϳ5���vU�/��%<Q��I`�a�8*g3�UJ�YhV�~��BG����V䃏���v����z?��-M<Z<�O�z.�j�z��콂D�0T����G0���{H]:�ŷԧ ;,��k^7K��Af�wt�n}س�/y���W��CmXuw.�"�1�.�Y<!��"J�K��@�_�Ǐ�.Xx��M�mL��K����	������Ⲏ�{r4oeY�ѭzL˸��&'��]'�I� �BjD�!������0`�#���i��Ю(H.��C���aQz�HڱS��y�7��@�F���:�ȼ�l;bюR�U%?�A�6K��g<y�Y�}Ъa�����m�5�C¸�O(����{x� vWI��u2�~���(����{���K��]p�Cm~;���8{���Σ���x%�嬏)jo,��,��p#�ǻ�ľ9x�d�C����գYjp;��+����QwZ��6q�:\�R�p+�V9�a�gQ�1��p1S�~3ѽŠ�݊b@
�i�Dٗ9	�wgV��p������0�M���^.�n��W��B�D�:a%�ͽ�>���@���iȴp�[8K��3}��F�FE�(�TbP47N�(=,DGFj����r�KS��\0���=աL��"��n��Y���Ɇ(1����fm��A�l����V�,o��8V�����WV%��������ݖ���kBY�#�����D���%�g�� �GP�����i��%�����@(�fJ�ձU��h<`��)L�/SN�|N�Y�'c�)pJߊn/�&Z��y�T�Ў�B��i�!�է�I����L�oƉ'������HEGr���Nz�J�X�}���8���}�A�g0x�J�˫�@=� ����C�RrR���XV0�sX�ᗨ�|&�M�|��x�S�a^*<ֆ�h1=�bݺ�y��L[c��f[�I9��p��]�Դ���.i�y�9}�8?�h�Gg�n5R�RW�����pЭ���Eʰ;ǭ1�QZ*8� ���%Tk���e �5G��Gԛ����\��p\��i��)P�m��P~nzd��_T��$!�Sz������U����Xʓ䁈 T�_��6:�' Q\���w'�j��	q�g���K/¿>�7�-]������=� ���Y� ����W/��a�S��Ch�����/���yG
/M�ޓBI ,w�i�w}1k�;M�r��:���(���$�rCdW��g��ݫC�yG�� �0�!�\�lj����o.��obo�O/+�u��5�&�tTV]i�?[w��06�k��5���&TQй��OB��h�>*3��5u�����{��A��U�A��|}ÁO����hz7���ʔS	�8��M���&r��w�m��i~�̠s1s��߇�,v/F����o�iA�b�s��sh��^b0�rZ�p� 9������<���T�?�L�\���a�X���/��ޠ�le9E���E�F�\#�}%��V�)��]���FV�QN����d�=�y��ǣuBQ;��Җ�P��Gk�M$a�`)��/�Ro��"y%08(&MHM?��Δ��h�.�e�&R�5 �ɱGC��^�lq��;T�Ó�]�KFԞzC�d�]��uc=>��Nj�eZ�^Xx���0FaW��gė��7u�x1us���mоF^��?vbaNVT�l<��۵�nF�".��K>�e�Y�[v���wg�ᢇ�hE��U��ɇ{�J;[��fLI������Ӓ����:�V�����y�Wd!QG�BG�1:�c[x�g�
2T�ʯ�����*9�����I���e\}��N�x{��anuU�kE4����jmə�Ў�JL3Ω�����z�[����6���ḮX&|�&1q�S������R��9;����|�쌳��mF2t�$12�|s�sD�����q&�W�@�F�N�8����Y�%�m��.��Lc��*lRH�ܘ��R�T�F~��W����Qf�+\~v���~��>��wr��d�ؾ.In
�z�@/����Zu�1J��N����]�s1/�n�)�����>hy!F�i���X �um{wL�G�ʎė������IJjo��W� Bc/����[}���ga�@ܜn�>����6qY�:Ձ|/{Φ��aQbp<�c�m��1��lG�+]޵<?��u]����:(j1V;iJ��!%5Q���t���f�W��$W��������6�F8��[�%}�Rb��F�Hж����5.5��3�^���I������:��C��{���F��oM�XI�=2��9D*1Yݡ_m��Bo�c�ʀ5���v��Ո�T����k�\J�Y�D�;Zwx���v�d�����O���?�m@Eɤ������W�����D�XnM�퐃�����!�6�,�>���W�+Y�q

 �\��=��bP���CY���Y�.��AIH���65H}���3t��\��?<d�H�%b�):��b/w�o��> ���*�U`4�)y{n�<�B�x���͔ �������:d�_Lc��1]�"�;������x�C��Ƥ�`���ܯ�'3;(u�Z�,t�&�ɇa�.YEX�46�u���=q-�����-� i�8Y�"��o��\��L������t�&�/KN���X�2eƻ��Gp��l��y�
B�O�HH��<z�Km�j��wa�/r%��X'�u+�{Ϳ�J���U�I߂��'�[ � �E���f�
ϫ����c���	���K��|KQ���R�IKN,�y%���>ZՆ��$���X��\�j���'neP7�'!�@4���,�ڥUuz�"㱅���*ڠ�Y1���ׅ�np��_�ߘ	I"� ���޹e`���zV�R�OWW��ɝ�Q$8@�|l�/4����V�( ���7P�t�>R���q���
oAJ�N��VY�|r��\3֦ms��X7-9�Z,;�SI�U˹��5,�y�ۃģ_����)�&ђ1�����6J��r@-�pT�* W�l�#�E<�Y�+���J4��jfg���7�����Kx�y:E:��ɾ��=欇f�r��$�_�I:h�
8�qK�� ��Jzy`��"�s������5�-�u�L)9��Ս7�	¹�5K��PH��˫
�w_t���S�z�~���]�u��٫���BC��e���z�;z���C�)Uhq�IŻaf���$/]���z�E���7Tp>{Kf�M�x;�)S���9��%v�����J���pL��C���\<��6���m�4��~� K��A���1(�-x@ì���xL�k/�*��xL��n�|7�S�P����S���ݗ.�Z�[ָ4S{9�V�QR�(��;Q�����)�w���r�1���	=pM�SO&�:�]gTy�O:���o����SoɊ���ߺ\���|m���ݖY��BW�s/ڌ���Pj	s�l�=.	\�(]�u�1p[�	�\'#X{C��jJ���6ӧZB��w�%�����~ܙ���4g�W
L��Qb>�4�c[��
6��}���C�3�(��\�g�{&�=
?< )�o�!� "g¬KϷB�b}BE�D1�̌A���^U�-٧y�đ7b���5��9��feE���Kq]�H�EL��D�,�b�t(������9�w3/��<��2&�|�.,�Ɏ�����(^���`@�e�B��*ZD�)G�i�H	:-5�����N��~��P*%/1fk�0l��l�y����Y�p����$�s��Wg���(��������m���p�w�
%d����?[
�hE�<�N��Va���͌P(�;Q�Ĉ�˳�EV�ƣmX* �h���iӋ^��gB\��~�\PR�%Ԇ:)v������V6�������/�;Z�pZH��q��Y�$2�����'�tl+*ys��DY��  !��a�|��`�G���%R4 �[~��p3�1M8���}�a�M�bpD|y���E���|�H
��{�6���G:�Ł;���+�R�=x�`j#q�,�v��88-;(��A���+�v��n���&0_i%����5Z\�7�D���0n*oG�:6���"YC��p��͖��a�p43��`#����w�i�]�����~��]?�F�f�)b����f�
9�sN��*���c]=��K� �,\-:�gJt�_������$�
�5n���V����ق���!z�լ�p]~�
]%�2����M)����7\��e�U*��Ow�:��6eKC�cu�tK�l��F�Kj���2P�M��7��b��q���/�����p�:���v��j�f�W�ĩ>f����$;�[����0�H��l^�J���ve.�\�h�� M_�
镤=�)�]�n�|d�^��gçA��"!?nAt�n#�P�xk�_�e+��^FϨ��	sl��91)�&3њ����W@�;�qfӔx�S.�u쭲�eu>@�(�LlÓ[�v�.ډ+��Oߜ�E���E9�#?��@�E����>��|T		��j%ѡ��7+���-�(1����H�+j����z:f�M���@����ȲK0����Pf��ie:����m�Y�Z��]=3�G��'��{
���I�"������Qd�U!5o-�mcd�c�!x5�'��H�\qlJ�uDU�*�Y�M�������zbM3/� y�1�(��)4��s��Yr�7`�S��ס]gL+��H8�d�j�(�:u	aC�)�}�Vv\dp�g�~m�7�Kx�B�4	�Y�	��V:%��,{=�1�+���'�G���12_|BUu�D8C���������h~����#��Ll��(C62�.���u߷m)CF��+����Ne1��� =&i.-��"\���U���S���e���r=�������3@KR���}���q�OE��;�a��k�f �G����r����vR���K�wZ����"�'�EX��+0��Xu��csnQm�췣55wi|��SY~Y6W����wNi�xX�#���f�t��*Ds�e�!l)"�~%p��c����N���a�i��GXɶ��v	Uy��Ǔ�z#�9l۔�W�������ɉ�#�Zt�(��j��^�4!�cpk�UyyLO"�Ys.����ʌ_4�F��Q~����t"�|�W΋3���;)|p��쁭�?4"�����8X�3��Y����ӈ7�����ђ���ˬ;�X��i�%X(�G%֥�RV�P�9���s꾆i2����c @��)�DkXH����
0
��aڕY ��t�U��쨅QÆ��V���w(Dhv�m��n���<ճ��l��.F���oĔ�:��w޵�H.N���&D����ZE;��S~�H�l�(�}va;���)P츎��j���kM���z S zu!ݜ��&�V�DAa�����w�!\'�	˶uC�DRw=F�Mj�Z\;ɐ���ŉ�9�ѯ
� �//[����| �&�sTM�KMSҺ����w����?�ubB}�^,�i0��h2�h�̇a�aV��������[�U�NQ�� �f��K�h���f�ԧ�y�'�hB^a�2�@��Щ��t����_S�ӆ4��(ЏP�\
���A��Hb�'�Z&z�`�3��N�s7忐jl/c���҇K"��)k��_�o��:���I�(9:N�Y�\�I�Jy��gK���{���;��ōr�]�z�����!	��q�)pi�\[��>�rnkͤ&�f>㰢>C��Hg ڥ.�7�:KAf�j�p���)Y��#�"��fz%c>����M�P��
Ud�?LUf���(B�H��+Z�S���Y�`k8�|��->�ZVw��o�Kq��ӛ-1̆�䅮�6f��EI��
Q�jev����@^�7>�#~�җ���M��k>hita�@6�5�duޣ��'�q�X������z����Wډ]#�[���2�OI�$֎�?�V����KD��꤁ψQ�W�;��v�p�ּ�o�|�_�j���R�3Ãv��"o�U=�V�L�)1 V���`Ȼ�m����'��=���p���l������~%>��|�eغ	�>V��S�9�a�>e���+iv�T�"�)�H3;��ԃ���U	EQq�CC�&g�Z�ѱADT���$�[�v�V��d�_c�
[��7f���t\��C�ث8�#E�jg6��`�^����R�+1�ʐ����6īc��,uHP��_H��`D�0F:�����.���e]+�Rq
4.|(��|�X�JL�8�:������ƙ�po���\���77�*�]wByu,��M�9Ȳ	(�C�d���zZ ���PR����g��C��yg��\�Ω���p�'�f$Z���	��d!�����n���6��u�ga���� ���.��-h�M��y7�l�lyj������}ӡ�X��cB�J��{ 9��9�Ka��A1r.�  �ê�_U�s��n���3/j�˗�x��ٯ(�*���6�ںj�1�C��̮7N�*����B�f$���ܼ��`L~XD�=�C
�#�B��=*�"��H�4���>'L���)KRGi�zX��#<΄���x��bLH�sv�JE� "!B ��c�_�AP���%2���^򖱣�G���o9�?o`lEN�b������UA�ɹEw��k7��i��(��d#}!�׌�oR$Ӭ���(Ք�{Z��w���)>�ͬ��7��8&(�T׼{I�oi��xn�vM~J@4di�V�K��[u�1�v)�pb0�K��m�E�&%����0����̫�����?-n���;�ί?�m�>��ʹ�8�MG ���7?�oa9��Ԋ=������|�x- ��E�C���ѧ�G�����`/�)�����'Ot�ҸʷPĮF������x�>҆ޖSۇ�a�H����K�^��˦�o���8�6�5|
��	�P<�χ���������,�;��350�㞃�0�㷨�z����rID�|�ٯ�.��>��0�ewY=�Sc���vP&a�Ƹ�ጆ��*�s���#8�s__��2�bd��- �b��N�=AQ�
�xH�d|tBu R�d2��X��Z�c���u�b��ݶ\�a�d^hC
4؁��\�"�S �]�6%��w� �(�'7����Ә�ŕ*��D=D��^�;��� L���c�T豄���9U.�f���iߘ\�J��ԛ�	�RG+h)�
㨓PWR5`��}���aBl8B$ި0�8z�����81�_�(/���R%�����Os�"0(u�ч���9���!��ĕ�9y�̚���rL8z�AQ�٢��
_�����(:hQ(f�Z���!�23���~�q���G#yUb�U
wdģ��I�\����E]J�����A�CD�f��9���Z:Y�o2�!sI�wZ@;O�p6k�8=�z��49�p��s+���l�C��q�iEI���J���q@A_����m���A�H^���qI?�x� 3��F�@>��^�0M�!��\�G����0��ze��/#F�}ak4�X4x��ǽy$�BO��"�Jf:�~O�<`Ig٦���(<��n��UH�B��f,��k��T���#Ɖ�1j/|��6_	+�}�u2�+Ǽ��~��<��0�b��%�NIھ =e����i]K�\��غ�5*�S`@����߸d˞>B���
FtC]]9�Q�M|`I7LRK��q�IK�l��U�!�eA�ٔ�ѯ���=f�7�I�(�r��YQ�ǭ<��� �qE���)�zJU���U� �r5�|�r�ma�(R&�Fң�
%Z���,��#)6L!=ܛ�3C.�G+IF/�pƉv�z�V��C%e�g,u��~$�
�z����EgU��ur�q�1��Sձ�ߗ�5F%
.b��yQ�XO	�av(׻��yan�n[l<�\@}���
-��엋.XC�}<�h���"y�3��r��gڌ8��N)�3��#��}��6B�u'4p\ ]�_��4�#�@d%΂�gp�Ie����G�Ñ�L�Ͳ�����A��,=t�.J?��J��}�VjA�lM~3�u]o��I"")<�4}�Ϳ�iBuu�S�nK��9�����5A�[��L`FO2��}�]�p)�ہ�u�!ĩ�<����ՠ͉̳�Mv�������-��(���.�^��q>�������������U�����qW�`u�L���7�s �hS57�Y���������r�B��7z�lpZ���*��Q��ϫyv�v����@c�֋��ا�q��U��ƅ���'4mXN�B/4vao����	̔ho�U&W��H�*�����e}q���� �����T-�Ƃ��w��L�+����E0vZC����P��QIBxH�P�ƪ�$7ӵ��W�^x�C��P��/����M>�;�h~5�(U~"��sJ�ئQ��o�۴�m�/�o�vH4��o��Lģٹtb���ʔ4��j���B!�)�g���ߣh�bRBѪ�C �شd�y}*��1�����`�s��	�0���I���+�N�`��:*y�xl��Q6��цc��NԞY<<<%�-���[r��	d�S折��I[V��l�L��~6U-��bqT	>)F(=;��ӓT [�����6�:���D:�m��d����_!R':ej��i'Jw�T����Y��w?�r�p��z����Q��
_c��Y�k?a;�k��֯)7��n��!��z�O�ׯ���6�1󟤓t;Z���}_?�W&J����|�h[5W�#���a4+L<��A�Eb	w'�AT�𕂧�X��0[��߁hw�HokФ$���(5?�T0)��>�g��]鑶��߃�9�j�t�R�!Q��/`�����S@�]�'1q�%%�ć���NJ�.���2�DLƚIy���:4�wĺ���#�󴨠Ǯ .mDWy�3�����bAE5�O�/G�O��<[$�j��1��tg�m�0k��	���iVѓ���&ch ��*�J��ow�����Q*��j<��L�T�=Q�=�e������gAۚɹH��Gs�@��g-�|�A����V�E���&3�B>E��z-
�z����𕁴�h�Q�I��s���YȯZ��Z��a���G۽�:Z���|il�b��**�ve�GJ�+�8`����B�F�醄�׶��w)�i��� �#�)#R�6aZ�F�f�� d��(�ֆ����������j�N�;@a�����)"��!��8�+�|p.؎�NN�������绔�6� �;e���P�E���K!K[��B@`u��M:�2Uʔ��[ڦ,�w4�vq�Q�ݼ=Q|��X2f��;h]�K<�^7�W ��*4T�E���0�����j~�g��Q���s�X0k�W��wda����Ө�b�H��s��W[Ɩ�ڶ��K/�K�B�����r5���&p+�q�4���˦Wl��y����e��:X�_(�ZV��I��ӈ' 4��Wei�<5� g���S0���D�JP�Ly@�;�ϔ2y|�Y'�!0�q�|^%W^�lo��\��/\7lN�Т�~5j+������P�R��!h�-��{��nMV��O�12� �Q]�^M�>g)��v����n�;�'E�4�ケ�sy��e�>x�/�
E�=�B������@���ZC�iY�S"XO+mB��z��R��Ln��e�H1@�[o��:��ïfU"�,�_Ya��3���R�g��_�XK�R���i�;�����*?A��@YM"0,3�Ki�a�99�,^�*=M^��S�x�2bc�[\�&C2�,�
[�\;�'�Y`��u�-��-�a%I��b�ԙ������ڵ5h oFXL&(�o_��X:)��l/�@k��Z��a'D]�8)G!1��$K�u�X�D�����n�8��&}�Dd��+�l�3i5��f��%��Q<�B��EC���P8�֛�גo�7>���,���-��6�uq�@W>���4)>�~����;�Z"z��<����A�8����@Q�
��&�}u>����x
��Ix1qR��Y�ʅ�E��C�Z-�Rtf��w��Y�'8��W�׹�oѪ�#�2��T���X�i�"}���*d�%��d����u�9Ҋ�i&	$-Zyc��7�2�I�m������|�!,�u��Q�0-c	����c~�D�.v������yx��3��|1��%'<H� vV#�SY�3�dG72(A��ԉ���a4
H�$�k�D�fb��+s�jW1e�	�G\P�ab����eM�^6�P0F�j�h,֓��{�M��$xp_8bB!΄�O"i��u\���I�-X�X)��0�Y$�$���h��0�z�"��	e�#L84��Z^�
7���-9�� �2.���F�
D�Ψ��K={�k�@�=�����0	H$%�iK�_�P�Q5rw��O�!c��eO2�)���LZ.<c��;�Ђ�b;����0��/�um�˧Q�Q�Е��-n\���7X}�,���#/Σ��i���aM��/�*N�t�r傄��x��k!5ȉJ��P�ZCs���;���R����'����	�:�O��:��6����<����}XW�����DtX��Ns���_�?��B��&�F�L�[�����%lB���;E�&��@;۾Ͳ�����K���j~2�%���:�rW#Y�G`D���rvqx�lA,����>�,��Q��*Ή l��2K��"p������p+#�֍�	�)#����çBL�3���	�;D�99&XJ��F�y6��f"�w2�r����xD@��A+�B1��Y �agرz�#�3I��#q�ވ�+��>�Qo �@{��4���qၾv!f?_Ӈ����\Q���z@z�����V7�ׇ��|9*$�YO��:��/mk1�d��v/�W4x��g�`�!$M�4~������,����z����h~��?��Q�����S��,�0m�g<|ė�q���5��)������\n羆p�g�!F�"�zP%�vO\��8vQ�RC�*(z���V��~8�E�_�+	��繛H��8�M�9L�����4]��l����?ī���X6��*r�V��75�xwCaS6PἾSf��g��$�����Tٔ�+k8`��su�$�1�@�91���$6&���=��Os&!�or��"�
�,N��d)�w��)��-�-&�wVK���d�d�SF���5�t�C����]0���Lpe\�(y)}�1��)�� �.�.�i
�`���`��Ȁ�R���Ɋw�́�@MNK
��fcdi% 6��z�Ȳr��Y���*Ǫ���7dV8#bo����÷L�U��e��zS?x�����݃��4�I�?��DE�k�ߓFV�i�j�}5.y�ڣ����_��/]o�x��mF�`�]����0Se]c��y-�"*U���g���m+J�|�&k|NE\:.1��CH�q�Hh���VS�KZ�%
�\m,��%��lA��T��RY�"�#��)X��n��]sЯn��[O��kg�](��O�f>��e�:e�u��i���t����l�.C�1������E��ޛ=]��=[��,:K ��ɨ]�Mo^�` N]�!L�9zX��fw��I�R�'��ۯ^����\F���� C�Y=���*-+u��~�n���9�i9F�+�Wh�F;�68��y.�3l�T���p�ae���9m�P�ؚy��h[<���v����ՠ-B���wAd�`�����!MGl������7�������+C�P���q�K����ۚ�����IB�]ܔx��2�(�|ù/	�%��|P�T]9Ӭz��n-���1پ?b	e�x���|E�#�Ӗ���B��dhi"z.�{�~u��E.�!�?[�f���iMj1ْtB:�̃B��:� �y6�t���?sP.%�}�s�l��j�M[Ɩ�,Pm-�h���|j0����sj�M!گs")���'��3���������E�"`4��t4e4�bT>������E�U���/�}A���*o2wZ��z����g�|d-d����oڊ!����0�a��!��
��{�}�C���sY��^�G��䈝1̷�������9����o���$kƚ�,�{4���7pf^�� KD�Ss�U����#�o�Ɏ�ېQ���ٜBǵ}�KɊj�W���g�E���wNB���ʀ4XN}��m����&@
�i��Ü:��.4���v�א��,r�~(X��рl˃t���>����:d�"����`�-)V���x�$G����|v��~AW\�5�f`3��c(r٣�Ӿz��1Z\�����ڞ� ܎}xG<S�&Y��������=��Q$@������8�`�q~HLaz��H���3�Y�B��~�J�.E�`C��yH^�܋�Bi�A���pm,�9����3����ٹ$�$x�}1t�)Kʅ)G*��"a����G�_�V0ֱO�ʟ^Qor���9�����"[�ZG~o^,�^���Z@) �9����NA*1~�,��[h3�Rvw����Ӧ({�#�W��Y~�y���?>���iZ� C)�Rz�ivV��ܓY���N�22���8��Zũw?�x엉Иv��:.%��J�O2!9�@�RL�0v8^�&�h&�1��Xk����}��!cJ�-Q�'��_o�hu�9
ʫݠJքq�/C�
⬻ׁT�gNU��dl=�����e8��5�Bl�C���LI�w���q ��BpɈi������K��<��ID���©Q|���|ߨ�&j<s���Q��C�ja3T~�!o[�Y��Y;f�lfJ�;�z�v,��t��Ay�y��j��h���ʦS"/Pҏ�.�=-�5�{ >Uw���V��lIP�["B�V!���t�@%�Be�1 �d���8��d9I�e�Zh�/���,��nqu2����> d�YP^��I#�]����@+���E�N�oͰ%]�%������)!�$^Ec��a��3OlwQT�������;�k������G���ْ�`1�Iӽ��R�/տM�,��q(`g�m�Bq�ȡ�D�MPok`����Ĩª��>��'�F����9�h�$���^�^>��	�y_e5�&"���$*�͕%F�|����_7��Uv�0�PǊ[���d4���G�O���z��}�Y�'cXLٛ����ŋM#F�7�,E�%6t�u��P�a���ծ�c6ڶ �g��;��cϿ���u!<Ek?� ȃz�-��x��X���5��қ�9{b�Ef_��J�޳�q߱��L]����K	V�q�u3g���RF���-�)"l��P���޵捌��Y�i���Gy��o��;ʶ�7��4&I�x;1��v��;U� `���,�BpDpڮL��$�R���{����+��v�L{Y=���'�hA�Ot�#m��ٯ'�h�E��X�_$����q�[s��י�1%�J�`j^�� w�Ã�&ξ�d�f[�S�)��k�ѡ�=��u�E�l+qS�}X;ti3��4���R���;Jx�L��׆)Q<�Q�h9p8�Vv=m���!˅Y�؀Tm)��m�.
��`�:t�Cm����3�7�=h{=Aw���L5kb�A��V_�M"ƴ�u"nGf4Ŭ�Cv�\�N�_�����L���M��4j�f}eFB��}j�.I�Hܽ����M����lV��e��Dn�ٙH��/����Ѩ��G�%�6��Q��p�{F�o�{�����2�N-|�Zޣ�,�Dŉ�zۍhQ�.��Ĵ�����(*>U݃`Ӑ��Y�+���%���t��8Ayຽ���N�R��Cl�< i��o���ۣ8a���5P�_��ꗞX�x�M�ą�M����{�tk����Д+�Bm����6ʀ:�)n�l´��������A��\H�Ć؟�2<�plw���D�f!3J)�Զ�^�<�W��"U�����U�@2��EW�Z��;<~�S���D��>�E}#o@���g#$����Nܾ�c�%	��z�x���꽓���'��I�� �X��XM�L5�VXl�T�hk�Y�9��&MO0�^,��4O]EA%���&:� ((�e#ӹ���;��R�u���z�l8�ȼ̯��P�k�����~Y�BP�ے�sV��ov���:O/� ���+�'���5�T�d�C���g"����\�������
3�C��L����N�=�(m�vu����y���bo٫"�_�=J�`��� �0'��ȣ����µ���]���!$1;$�J8O	�ط�h]S�dfdr�\E���9+ߑ���3�77�,�{ߜ܉�l&�=0��@y�/�&D�2
n�ќ�F��\�NMഘ���m��8�P8���s��E-D�9�y���o�S0�M����5U�=��(�ҏ�,��Cx��p�>G�2���m��ܗ������gI��L�U�D���������rZ�fv�R[D�D)�]<4G�n�پV�A�_��P���/���v:_7m�D��r��,�4B1?+����e.��o�Y����+bQ��>�[3B\=�,��ՆY���۞틉V*܈m)��4E	��'�����&���)���	��I��F%X�� ��}b�GWA��0/��I1n�4,w|"x�&nM=ԝ���h����1>�Xɧ�h�&}��6���1n!�3���&'��g92�}������d.�a�a5��ǜѪt�;X��+g���%oh���9?���ɸ�Z7�΁���G���_J?�k�H��]1`�/�����T>���_��8�!���ݺ=�x��D.���du�7ǵ9�M��%!�a�����csvj�+>�ƃS�<=QB��TF�▔��oӪ_���I��'��#�%	�ldZ.`�Z�Փϧb�uEXin�o��R��.�4�N�z�����Z�6ܞ���ʲ����*e�f��UI��Y�&�k����R����j80l���g�!��zTbF�X�C��,{�sgydh� M�O�5DK]���R}��<9���8dj7�J@�16�C5v�,Uz'q�j%�H����ډ�d����|�H�x�k.������X����~�Mqr�^Խ!k�v��VL��i)o��<�������=H�j���{�M�{�Cl�49���xKQ,��'P����h����>M���?����cJT;����(�W����[$�z�s��ܒ;��O9qɢ�@)����L����3����~}�=O�@Y��6y���:E�A�g����[���C��;��jB�c,W�N����I��@�=��n'���I��v�����V�c� ~gxA�|�m~h�cZ��npʕ�����(��z�s2Nr�.�U�m������ȿ�/�6	+����^rx��#bo�k��h��(9��@[�,���Wl�BA�b���]����5¬�m', �{i:�َ�t��[5��* LQ�e'q�d��й�ev{�7Ӭt�A��ݱ�cq��Z5{-��gZh����b��>�h��?��j���e��HC
�zS<���!D�-���_8�# ����Y���N�7m:E}��X�v�%�\
�'���}�XN�bl�n��h��ܿ�4C��}��v���
x��T��MX-Ы#��2���#�0+���ǩ8EP~����p���'s�����N5~�VF��G��I��u,-�2�E4��@��Ԓ��;��t��5��3�����Fuީ8�kB�`%W,�Ŭ
����p������^�FKH^K��`��ѩrc𽥫�ըž�!�a�=%�5n���6�#\M5W�0q|��<Z����l�u�z-��}PDc��#qs��soZ[g6�f���Oq�A�OE�����ƏԎ����0L()�*����t@����Kqx�V2�M:��1�D�Ng��,5T>'���`���̸�ϲ��{_�[{������D��P��fv����ZU5��d\��=e��_aGi�\�{��w �����&�9���d8pE��R�$.��Lǰ�-�WB�1�*�����s�ؕB�!�w[��kt�!��'�̉Q)��u/V�Ն�8^�1���J�	��	������n�5���M/~�F�>��'C�.�� ��S+ SشAĈ/JR"���1�|J_�l9.F|���c�9DZ�Ǜ`��<�_P��}�&�KԡnW]�uМ��`̰������#����jXk��嵲�-+h��YGM���m��HA�-Y5�V�e}�$;!?5���:T'D���]9�o��a�}�m�^�?�cU�|ᅀ6��x��ȼm 7{��"��T&��z+�Y�.ͨ):K�-e��%5������`�p�-���ߨ��s�W���3V������}j;=#<��u	W������u�w�����0�@L�Pe�N�v���O7��r����q����&2�Q�n��*bG�O�.���d Q ��0A\�,觃uZVy'KZ�T"��Q����ɱ���!`��Eq�z��eFN��� �ch���_�a�ۺ�(~f�^U\���yT_�󌏐>A���\b�V, ������pc�u��U�C�#�ٰ��Q/L������P�+d#b~O�E���o<_9�)/՚�<��S�|@��z��1q��՚��|��<bF�u+im8���������ޛO�T��X[I@Y���|e�����"I��89�4u%��Uc�����QGWY[�J��Y(:X��Fe[��tJ��ჄG���; -.)�_�o���G�^{�����$;u&�Ė�f�dL��[�\c�"D��j^���ri6�&z���5�J��@B"=G&����n��M6�قI�v������V����#h�J�z�n��P�9�ZB�2Up'���վ�IAR��l���C/J�λ�k�M������ϥ�z�*���/ȋ*1@���OW�q����VZ���ԯ�p
2��  .F���s��A�����Pv.@�p'�}���.|���f4'�	���-�{�$2�j����撊��BCbA��7�w������'M�E!����N|�Xk��r�W]�Ix�v�b{��;$WŶ��ӝ��>�x*��p^�b�mj~���'V�1]k�Ι>._�.~��-��d$�$T@6�k��F���Ӯo�<m1HHk�y���TQΥ�+p`���*���� 笳��6�#��*f�>�zI5wT����>��J��h~��t�p�j���
ܠ�ZW�q�m�8hj�i�M�
$8��0��+9!�N\��d]�t�E��9���0I�����^���͉q(�n<~7p�(���7��u$�4��W<JĬ$��j�9݁Ʒi��6ïfI��1$�X`�~�s��y� p"���4_��x ��Z�qF/~S�M�LT�"`m����ls?��������*��'D��_YէW  
�:�g�[�zp&�PW~���݆�oC�˫���iF���gx^��@�ן�'��Bi�7fK	{?��d��D��r�j��p���Q�����������j�41'I>�@x5cL���ouNL��e�@Y�,x׶훔���
��r�/*�M�h���S�7��֗t�j�uv>���f�l_�v�08��I%@c�	��,������%|�Hw}��x;�����ջp���P��ߦ+���Mw�!SMΒ�2���|�y��)[�v������.����V~n����k�1����ԧ@D����1x�C�`D�[x'vq.]u���m���L/S���%o�zGyZ�E��p˱�����{9���U�����R��a�C���IÈ��B�����/��Y��n{�Զ?&G�x�ch1_١bDlKʭ�����|�ox^���Hkֳn@`P��2�3�������RF�=�9OIޏ1z���I ۞@� i᫾�s�]��c�h*�vF�����p1H,�'����>
��!��V���|��p�!��^��
*��yS���4�:���.��)�ؘ��z*�"�?d��v�l�H��b������Y��I���ݽY#=�Ww?��/-8�م<�5��#*t�f����S�4fuN-!J]�Q�Z�Pl�~+~,�����R��|�}NWUi��5�N5�x���DW ^WJ �N<F�v�����9�Amg��ܶY)���sZj�� &M������TM�L���p����^�G�Z*�J-���6���[���	]"�}�#�t�E�%BH�m8K��E$r[!�"Ť�n�x;	1��nX�_X�okP"��p)�0
���^�of�^��e�HZ�Ӷ��Oct�s�#�16��&<O���ɥ� 9��,�3S2�l���D`l���x#e�<�2ȍ�C�+����.�c@�Y
��h؀5�VJ��=
��,n�*�sf������k��ǎ����F�m���,�݋�����!�&�h {v_=�l's�,ǟK��:&��$m9kW���e=�R�U�x���Y�-�a�[5-\ۆe�S��4ֽD.��Y�V�5�2�~i}��(\�"�͊�s0D�׉����<S��q3[�Jw=�ez�B5ct��Q[1"c�#�_� ��b�������$�E���9����5�h]fY��(��XT��kQ�ޝ�� ����_�yo:���i��җ�q�*�y�U���Ckő��4F�
&
�ZyUT�������~���cmb��~!-��:��4��1J	aسP��V2���%�]�����<���k�<��@R�?���607��δ�`d�0�;���eT�a����`P$�w�|�X|;����T��юh\���U�*�X�D�-FP�������p� �u`�vEW�/(6��G��P�,;��Ҡ���O��B��H ��;%ԱE���~�t���W
l.e�'��X�fվ�ђwr���j�3�{��B��7��bC�v�w�چ��7�&]b����h�<jy�&&���:&����L��6��48��7J����e �!�l/V\��_�!_��ӯfZ��.���h>h�cAP�C��F�����g�T��GVP��)z����q�b}4ZNM(~�	Yc.P��������&>�
� �<�L���u����^	Lm���}k�N���f�l5�F>,�����4�Mtm�I��9�KӅ��23y����7ۍ�f�Y�Xļ�2��})�����9J�؈�@���m��ٻ�p��t#j�1R�,�0�'����oC=�T�e(^�I髉x{<��&�rx�S�	�Hn�{��5"$}8�/�秈�&v�\^�ST����6�}���+a�C��߱42`P��PSxZ�H��N�PNaj*pC\��FБ�JH�ж�3��C4y�3z��L���ԗd�)�h�c�o�NǜL�9���k~�G�F������,�����iJ�ӎh ,:���:4)���O	���-R][g�4�.��d��>�C\W9Q�ʝk��V��-���┯��~����O�	�jѯ�G��X.�� ��o*�8�)@��tD!�\a�>#vW¦;�>����vlc��4x�Qo./����̺U�E$��	���`�e�H��Ϝ>r�czjȲ�B�`�=`b������%�q F��I��!z�	ɝ�V^@�)�Tm�̍n]�Q�\���ѩ]-�����w�����G����RPm����	+/P<Uƃ��B=�P@������*�:���N�,��R��<]=y��Hr�P�{��(e��ۡ�si([�[���-�/���Q��_ȇ�e!�j��Ʃ=�f�jo�zQ����3�<�+�$�o�ܸl8W.���'|�Z$7� +�qÔ�3�2�w.�Z�EK)�(�Zß�Aڛ�P�mG�RWO�K�>YkL���q���%6�*h� �NF�cM����NAc�������4��f�q� )nu����?hs۲��[��6E�K�or����[��y[�Lϣ�98r��Ӥ��1��pD%����U��p�=�ru"�c���Z��_H]�f�3��t�'T���N����N�#��a��K��<�?�S�^� �P�����1}!�t\HH0��3��<uz0������ːCG0x�e�?��r)~a��/S��� :2�7A�U�<����jN�my���\�ϝpa��p��ǐ�������[XI^ܙ6!�>��};�m�de�'hs���Z]o8/��	b�U��,�~�o{d3T��M�LSm8��|D�9a���K!��'��c
V��'��h���@C	"�������<3���e��~'u��#.��������4�:@YɗPB�vj��l%6a&.�S(�W�Ljxz�5�D���L�*p'K%N~s(�_`�|�v��Iwn|0��(V�����J77L^;�`qE�u^����f����fS=���mF��F5h�����ó
V�T��k���%���o�����]y�G�I����=M���Dq�2K�V�8o��:U�赳������zA�4Ј�4��.6�����+Ȉ�t���!D�R6evw"��cJ�-�������Q���\����5���u�9b���ɏ}��/�����LP �Nj5���#�G�:}}�!��q�����ZR/�u�,�Z�i���t�ö��b��p4/����(r�'F�U�fm��h���34@���l��G��I#>F� �����=
m��d$KR�,P�m��\�����d_2�{k�V����6u� �H�qWxo����;;L��6	�����ǒ��������F�A{TU���Ӻ���0J��QH�-���%=�Z��]*\ǝD�R�aҥCٲ ������[��{I��}S��Z����F��T�&�v��HV�ѻ��or��Th����ѳ�<���oA�2%�b1�%Y���~���'����f�pX΁ɬy
CF�-5�M�[�F��`����r�ߚ���aG�r�n�zpĢ$[Yc��}V*����%F�(���f9�����G����^_��`T<�6=��d�A3���˴��]�,4!��@��S�
��^� A~�pj��
F��'��.!��iT�^������3=�*�^O|Q�C��ې��`WO�!�H<��U��3#w�d8�KG2��=��-�����C�`���d�u��|('}��%���Q�^��9�~��
�dFP���8w���[�$N@����^2�I��>�5@��a|�X&MZ�KAf4�0�vHxw��]dʼm�.�'�!j��4��U�e����n��+u;$��&��%�����!�DC�� (�K_���λ�^)/�{_^�=�V��2�0�����R=�!��F�4�)x�[�*s�iO]�OQ
�@f}r�@9��/�ʼp�X��NP�wm�S�T��ޭ���!�hi���*	��3A9����gc֭o���Rl��E�X���_*���i7m�&�
��(��b�Ei�"��m����Z�S�GѢap�3<�l"��oq�i6�s��W!oy�M�_+�P��_��&��g�,����6@ ��p��!��^d�ALJ6���/מsWZ�ʒGh�GOJks-�'1�_A����f�|$�S��zb5����rg"	����N���S!8O~2�N���^$go���][���r�6�_�;8�����"�2`�,�)�;�9X�w��T#�~���	��#�"���4�B7���w	��W��jA���}^�B��M�%F��c�u{(5R��3ۛS���G��,.����S�`A���ֶO�����gИ���u=��vV� �����j�Ĳkg�i1���T����6gpK�Է�0�]R���IӔ���|�%7(�<U�K�駉3�3���� V23�?�:2E��'$*
��A_��xPE#��=?v�?�3�٤���M!A�C�&�g�a|�* ��i�Zd�\�Z
<������[_�s��`!%�^�|��*�]i8q�	`*]'bhu���<�n�2��5�	����K5��-���o/�Μ�5��:��{�Tc�cr+n%��a�c#.��9E�WgBd���ܼj��sz�#�����Rq$�Ѣ]Đ�}�3�i]*��5g%�K����ޗ"ko=cQ�i��@b�bj��s�y*�d0w�]���ӱ�.k�ܳ�i�3���2MT��>[f��Sol��V���Ų%��j�;�v�EC�F�I7Z0�B��#Z��.�;�Y��=�L E����\�@ф����[�5� �մ��}ca_n��p�V$�����Ӟ6͗�M��j	`}��DיAI1S�Lޔ�?��e�챜j�Mف>�G"�nK�V("*BO`�p��j�q�K	q�~�>f��u���fa���F��q��p_W�*�LS���������4�m��r|Q���;r������74V��$���[;����tr�i���c�Z�HML�*�O3�cv�	�W�P�oc$asAt�x�BW�]�a���!Ľ�f�B����D�_�(sA��8�1�>���%�qla��TϚ�"�-͆CӢ)U�M�G)���#�x&x��2�P����k)�%�'�w9�\���A�~��hnd�:~?�Z�ʎ��A�`�?B'�
�B����O'Î�[E03�5�l���C�� �F�ښY]�"�Is�}�J@_1�v������#��� �N(zK=V^5q]^��E��`I���B�#��י/�6Q��u]J"�^8��a����/.���N@���HP�6ēY^gKc6���5Sl�	���;��С�?ժ5����w�H&<�N+r�C�D�q�G�}P|R�h��v�Z��_��K����k�l ��<�M"�����~K�{+<3P.��ҥ�~<)z��H��ę�A�o��\�}�\��P1:H;�#a�o������N�BIK��p�`huIx.�� �Ț��x��|�б��.�\Z�c�Q) ��`�{��y�H�U,/�/ճCY�� ���%�ۑ"��a�(���X�Km���R�1q�u��@ς��$H�q�^�H�+j>�uӵ�����W��R��a�Q�`l��X��S�r�駩
v�(�-� ΰo4+A���TgD�]�:F$4���v���.���#"`�~6�N���6aabt��[�R�D�6�� S0x�b��LWg��i�{k�,�����	=ř����Ϳ�����6��$�ή�r�������l�(�I.1�T�}�ԆC0�z$�!�'Z5C��4U�amd���ᕰ+� �;�gxg:99q��p�V�� n(9�	���NX�P��d17��	�L<��T3��-�5βpe<+�~�v�9:
C.YzG���%s,1�zu]�b2����$�8e�9a���[h��%v�-���gbȫT�������������:�0�\
ǂp�/C��ߛ��-�j����VM�i:5Y��U Dac��L����p����wL5|T��F���L�d� .,�(i�#���u/���=JG����y�ֆ$q@ԛ���;̩UU�'�����.�`9K+���xD�f��H�Z�I��b���=�������4Qb>��0��ڠ`��c��E÷'b�B���)=v�,���3 ���Q[ͅ���j���_�;-�����(�_ޤ�zeØ�Y�l)\��0�F`/��L�o�,4��� ��8�Q�)���7�����ܲ-�ЊO˘�#��-������d�j��E1u,3*���D���ˤ��9=<l����FC��9"�F�P)��=�S�n�I*.l��gNh�]��$��rJ����j�����!JIa�^�
4H� 2p7im(�w���X��ӯ�����(G~[!�#ow`�hZc��ګ	qK@�u�A�M�ݺZ�l`К�kP��Ɲ�?�}�������~���ȱ�O�Gc�@����~�@�4�M@�4�0�G�Ak-�zA�|�ޮ+�TMz1Z�K���qw?8ԑW�L3����]O���U���4�ͥՏ�0t��-���.�Xa�aI�u4�� ,(�@	?R�<���hAv��;�ZVR�]��"K f�����H�r� ��v)ܵ��b_X�H�7}��}v�:� |f�F�������bn��|wg�����1^�Q�aN�y9�:�\\e
T���D.��S=U��w�S�m�ՊE�g���|��O*��4����	Ks|������:R|�����^ �*���K��ej��r�u����0�����|;��'�,���iX��Eq`��ɜ�Py�E5����U�!��Yv}A{+����B�,�qΚ������zw��ˣbaZ�ȌcH<᧸�E�M��m��� ���:b�rb{�Ct^�\0N�SO�ή��hH�Z/�<�x��y&V��ӊ��%p�KLO@-�^����-�D��hϞ}��,&��I_������1�bAϹT0�L�a��Nоǘ��h��1k��m���)}��s�my���l��`\�Ւe���G�9]P���.h,v�����:~V=���Ҥ�I�\�N�3ӳosA'����Nҹh�z�ݭx������u�����ཊ<@&�z���:<]�����`�i��\�7�[���-��?�&! }�"]d�YP�>�MhH���=��J-E02i�������?�;������5�A�Q�1Y�0��#v�
���6��V�_ЋIuZ�Fk������X�ϻ��M��H��o�;Nj�I����@�� ��~���1�-���Ǘ"l��a�é7͞d]*�8yƢ6���&a�������1�	q�r���Ͷ���EZ��@OӐ_��X�
�l�F�y��,䓪9��7�����a�9Eʀm}Z�>q�0cF0~1�tX��铹��؇I��s��Уh�� �m��4=7������VAJ@-Բq��}=���{�GǤo:q;t���n9J��&-���(�X��m��%��X][�S�����~�-֤�um�~�	��m�JE���e��{�3観��u�3�jL��nPE���n��@���	5�� ����I�����
*�6�
?���&�Z�q� �m���c�UM\�ބ��}Hm��U�vpz�L��+�%��V�N�~?J	l�U�&پ����Z�K)"� -o���g�{gJ�7@��M���ܐT�]~���Q����r&Of"�	�}��v�(sls���ڷ:W�S�u�<;��fC/���(d��[���o���G-���?�s�o�,;Tl�U?�Q�:��RG��ڭ��(�}��\r���>�H��Rc��!L��̧�es��a�f$(��L�hPW)�������r��$��	�DǑ�fi����p�8"k��@���s�9ٕ�A�w`� ��M�Ѝp`ϛ��������o��7I��}��[�Ǧ^^=����eZ{���hΫM��]�4����sՋWg�ě�����#����Dq�@<�_ǰ9��@o�m窱
X���٧�fI����z[Z4~UV)4�۱1��Dt��bP�fd���wB�BPB�T�bՁ6
���i�����;i��L�d�6֌k�pEc�\�朚Vv��tW�8-�ή��')�B������	�������s��FBd<]�`e�O�� H�*Ln3_�s�c���1缥9�~Nj�c"qM?d(%:����� jw�X�w�΁�4�Tg1/���N�
2��-���Լ_��^M����$�zN ���GҪ珓G�����50z��m�3h���ڹN\#@L.�p8�6�f��'��q� ԕ����[�A� �D'�;������sF��χ�	-��� a��X��������N�+��ޖt�tSb���Ī�B��G��j��Hp@�����SkX��r7̰G����s"t���~�
�.��3%�=�M�2R�0��)���� �
E���`K�,��qIO[��vX���ٔ_¯�xM�7�/澝�K��`.#�3_�_�[��kuz��C��6 �e_�
�:0Rn�c[t���ʎ�%y��H��R��w<��yGJL��l�XνG��!�Ζ�m�+�U�$5���-/�������,~�ъ��ѭ���~Q�ѯ�Y�<Xh�M�(�.�!ȠK[�fx�v���>s/����h<�[��!�����c��Գ�1������ƭ9� ��r�h���\B� �hq���v��u2��*F:B��ZRG��k�I�!�u�'�o��ִ�k�E{e�Z���H��Q�7��4�1�&h�p6(���{����t��I�g`�;�8�(D�
�Z���ce#)L�H����u��G$�a�4�B�nn��&�b�2N������ē�*B�:�l�"��?�������9��P=(F���'�ʒŎ����2�����p����Fp6U�x�@�Bm���:��5���}����Z���r�����ލ���:7ؚn��;44�탔)g7��s���/����>�Դv�J)��
�>]���LQu����X��t^*9�;�����*^�ܲ�$ا��|� �1!a��Y�p:���l�����\�+�R�5�2F����}�_ɭ�)W���m�G:��UR����hr4�[�7�e^xs�;}˳�`�K�뮱�������Ũ�����Iz�'M�E�l��V�r�v�,�rgh�҉l��X�3<=�Q�1��:P�Ùt�l�c�n�|�K�����J'� dhx-1:х��X�<�����U`/���*����,<����V��wԩ��Vzw�J�b��SZ0�\��lk�)h�#}DI�8����-�������2��� �U<e@I�[���6I���렍�H �����'��2����<BK���^]EV��|
e �oh����:{b��x���c�Cׂ�S���ǎ=�Ui�$'p�Y{��6�:٘ۿN�����.8c�_v���Va5���뵯۷w��J0�_\4�� �"�g�%�N�Sj��#�+^銼��	��ѥ�1��&Dti5D �:��U��_ �p��^�bAa�d6�V�j���m���Mv��|�S-�����.�΁��i&��8��8YN��p�Q(��L��\\'02�	�j���1/�z�zxՋJ�g�_�"I�mj��T����ϣ�CP�^( Qy��+L3�&k[���]P��^U���QfAkH<�z!l\��=&sv)䜻����
h��	�Ň�����Q��=��$N�<^�I*
����C�KXE��z��L���D�"��	g���
�Twi�#H�/�MB�9'9jH�6@��j5���������J�F������:s�w���Ċ��\��D�G�7�2��-�����?.��-�g։B`&�+��V,�s�,�����5�F.�P��u����f8�w��g��Y�^-�E�ɰ-aգ����\:�T��S!�̲�!��]���M�LF/�5���T7�u1����*�_�����,M��b�F'n���	�zJdO�����̾�;��0��>���t/���̓]'��@�{a@��w�y�p[^~�۲�I�U�C�.�:����.�� ����5�+e�����R�z�`L�F�'�&�ߋ�Y�q�g�*$f8��L2ύ4���H�(�[&����Z�9���n2�xA}nCk;8���;��E�/<	��@&uZ��є.6l���K�{q7�-
�δ�r�_~S��$Io��f��DΣ��n�&￀��o����^�VJ�?V�#kB=S4��V�-��`j�6�ں��#��g]�1<��uU7�_�۬/��n>���+|�΂H�~�����<4����*���9����i{\�N�]�e4w�ZT����m�	�;U�m�!�{\����%�ā��_OF
�墶 �Zb�8}��%��/Z���z� Q`���(���F�3n�#[�"�VJ��V�M�W��>~_G�J��Ѭ~ �,}� 3�|9�/T<`�^+8oBN�A3�6�+l���'Dg��Ȩ�%�}���xP������J�VV7NCiV�A�A��v���*_�1�4�2���"1BLRu��x.��1�`x����m�9ȅ�?Iڴ��dx�:^�*�l�|������}�oP�RN%���n63Uz��FBo~��^��u����5%:��>�#����)?���5�]~��"5�#({.�~C�̽Q�QƲ)6�8z����B㨍��J9I����(���N�x�m��c<5	m"�ɟ��v�	�N�en�2�Z�8Q�����S���G"8�eD�~�,*�����	ZϬq�̳Q����'�D�Y+L��jAI��4�e=�=f��(,��R��2�M(<B)��*
-&"�QD��w-U���������G�c̽�ŝ�їRξ�����ղ�W�;<�j9<�
+W�&��.�T����	�΍`fM"G�
#���\�я"��ۗ�&bg����_:���῵E��i}��b��E�$,��@��I��DsG��i�ܥ����F�K[Bz��s�X����k4l#p����N�Z�ж�[?*k����O�}�*D�â��i!�^��uR���4u/,��8�#��q,�s=���x���÷YK�tOn%����tSH?+F�5���3��[mSv���dܘ,�o�ޅ��*]tҵD7�-�T�y���K����):|���Li�[�1�%�(�ғ�Y|f��ڔ�C*/������*G�F��n`�x�7˖��\�`��58\�P�A(w+����gV�GY.�V�
��p���}�9�K�������c���Y1�,_�7t�ƙ�B���]pQY퉼�Cz��Q��Z}���51�0v����<1I-�d\@��F��eQЉ;u�]�v~]u��2=�p���)Q��0�OؾcR��61L��@p�x�L��-u�6�ߣ�|c�����S+��#|�� �vj,� o��}+{�^��1K\�T�W9��$�f���W�n��M1��Tb��'��9���>��Fh�37\z�_"��;�`��/l�%�)p��G>�*�"-!�Wi}*���
�;�5*Ϗ2-YU�^&y�7���M��?�<�j��Arr��.�)9 c�Դ[L��8����7�B��F)�V�H�O���o��v����3�E�S�ׂ�wY��a�����΍[�=��е�Pu1���\#���pzA�3���C�{�u]�^3.���N��U�ˁ.'�A�"��x�4_��>w���3��k����Q��ި�g`��%��Ac�븇6�X��g�L͒<�,>�$v��)^}��Gbq�nmU&������i^���dN�����vĊl�Qt8��C�����N��x[S5�!i��b�̊�����J��/qi�_|���su$U�s�Q#u3�7��p�B�JN�s[�ꐤ]�1�u������T�P-��@����w�� ��&�ℤ>�]N�X��x^���"�Ӊ�v$�wjBȐ0�%�2	��ȁT�a�᠋�����ǳ�2_E��$�@.�R�{^�c�����n��,1F�&E��'����3�ݛfq�8�lg���eܘ?��u#�4���i�?�XƂ��W����t9��z�<_Gl����@?�/�7��s2�Y4'�_��P��'L�67Ǧ�u(4%����n�dEz5��̩ȩ*�? ��bӟ(��Fb���,��;��X΋&����MA��-��.�H���t�Ɓ')J���Ln���{�V��R#c=匀�,Mc��I�������YyO)�b�[�)���@��Ѥe�u��fK�=�����`��g�&��ܶ��B�Mw���w�~R���jڬ:����w7��������ϣ��w�i�/r��lN��֠��g?�������~G�iL$�Bjm[:���P�3��@x7��ώ�\V�L�_���)2OD�1�?�ߏ�.�iOh!��JeM��7���#��
�D]P�K�H��=��J�Gt��Ր�D2����M��B��;�sh�:`�)�>j�,?�WU�i�v���VWq�vU�v�ދ��@��	�*�e���f%{���t���"��q��YC��#B�z�Jք��}��(~����L6,*:�6���ڎ�.��ǖ�e�8�����]R�2m@l|!�f˷�;���>��$��s_���%%]�1��!H��9�� 1�A) �vϊ�{��s��Ť#U�a%{\4����e�����&a�/0������5Ұ�Ɩ�/xt�1ԋ���E��I�Ĉ��~�I/�i?�/r2er��B �A��V`}q�7�%�jh��6:~^�V���$\����c���f�%b,9�%�o	|�s����D[8��=~3��Ŕ�~�pkT�X�ș;���?͟'�Yb�vR@�]�~O����QT9�!j���/
�¹�.!��0V��9�/�x�.�L2IY!��M;�3�2�#�d�8c0��r�C�&����T�m�}ޔ踖"S}�z/g���f��"nj�T���(�N��D&�UMs��Vy���߱<�I!Ojc�c�B�t�3?��*�]��!�F.�╴uR�A�R]O�^%{�wC�H���)|L"/� a~%4�>D��ʸ�D���r����%���R�ȯ�顁[�V]�_>L����vB�Q� ��F�ɗJ�6UB,��s���GB��}�+cS]���8ȩ�y�t ���":��+�<A�֛`c�U�LΡ���1���6��<;=^���Yv�O<�&�f���6�܀_��1d�lJ���%���o�r�̜0�����6��D�f��5�/��7O*��:/���P�>�.J�S��z�����H�AN��ߘ�2��a[�:*���$�߆1j��U���z�gŊ"�;��6��)ݳ�$�Q�kY]�˺y����)�!Y�o;�++F��P���Oqw���I����6��b�"#��.D��q!@طǤ]�[b����R�pei��sȄ�㕰y����n*k8�Q�E�S̓�)��k�����FEU4uG�Y~ #߯�B�צ��C�)�&K��R*��[����v�bP����joLC ;��"�wt�*�Y���|�����9p��~C(���Ws�0Za�]*�ܚ�1���V�\���HG%�$����#��Je�:��c/�P�b������P[�Wch���p�ٶ4�?�\�[� ggLN�C�"+}L��L�if��u1�ۜ�h�)���=������c�yU�`ʫ����o�dT�"E��&o�M>�yw��1����-�4c�8��7
�ɗz(!~P�tm�U_rV$e�*b���Sx�[��u{�Ie݅i;;.�Zt�B�A�)Y <�\ߦ��{�K.����_v�2�]���W�g�9��?W���TL��2k%�J�i��F[kx�7ER���s�،�X�:��8�0�ˁ�`��GJn�(�b)������|��F���m����iC,���$�h����n��T��i�:�S̀)Jt.U�<�c�����,��7{��O�k=(��/��;�癩�D�Z0Y J��h�ҖaO#��3�%�Xk�[��a�	�>ݑ����"��)���'0�|C��j��ƞc���	F�bR�)Ŵ�P�ߣEx)�*�����si{��8�oږl�\2�[C�z�=oW�*�S�U0��X,wR��'3�#�P
>�XUv�Wl��뚈/���1D�,n�6B_��#9	��:�e���@����%n_�,l=*L�~�DT����+i��^}G�I�[��s����(8��-�Г��Ӊ� &�Rl����fbMbY�]Hs��L	H3iL�!#����g*�c�s����4˓[-t�U�=���B�3߿�V�W�Ś�R<qPy�̆n�i��'��$R��$s���h@
b?)���7�S��	��y�I��T��
>��1�T��x�<�L0e8�5���ǈi��,����O����L=\��_��ػx_�J'�{��j#-т�I2���HlYӴ,aM��xX�Nl���c�q�;o�H��i|��*o�H���ݣ);��Ky[��e�Ud���c+�`�)o�zJ�+��۲�t�b뭀F|U�׏�C ���4O��A�AI��^���77���kSXc�< U���޼���od�$�g[�{��P/? ;��I�&4-�!�ޤ�,��(`�

�{�o�Xѷ��/��;i�(RS�@��멃[��neNf���'xbJ��/�zh�䗺V�+�@ʃΏ'���xNS�*D	6mXG���ŇvU��x# J��Y�,��|E�k���|<QevRp׳�Z��Xiϔ^n�q=�Q��OU��7��7�AP����Oҫ
3��&���m�y@J92rO���BT��Z]*��%~���
G|�b����	��Ks!�Gҵ̣+���}�F㧶��o4t�bZ�D����n���x�C��ϣ�[�J�%�?�b�0�ѝnѾ�9a�(MsD�JK�QV�u�k���!2[Cf8�@�K*��IVi��&�����A1���@�y���`�M��V��_������cJ{�2�Ms[�g�g�1�m~�.�����>��/g�^@���M'4�[�������ExU4�[����\�^z&ڪ]s��ު����n������Mmb��(�@�����gK)r�4;���p��5@��~�.r��$w�45X�K��F?��^LMB�It�����ο�)��ʣ���OA����-��L*"�����\XK���Y`RnƑh�-4�|��ay�ۛO����c���R��5�m ��Bu�S
z1Ňn*�u��i)\���A�]@eF8e<���w	GQׇ��=�v@d��ٖL���NU��6����Y���,@�U��V�7��aɥ������~XA�I��HM(�ʼ�����6����h��rm��ȾU.P�PF
@�ELsY�2(@G���_!���z���A�7���������;���-���~�X�h��n���0��8�{ d��&?jf�D�E��w�W�1,��.�,}���M��&.�O�da�8f#�e���t>N���^iӂ�fz���o���?��KJ�Z��^U�T�P�)Aȳg�4g0(Q��O�r�׶��^�.���/��T���ǋ�P���D�&@��7��!��8GZN\��wd`泀R쑚O��`�C��:]�ta��X�b����$��Xr2Y��/��`��c���:�٬�а���pGTz������8+��~�Pj_��C9��˂K��������y	aK����[Xg�nZU&K½�w�f���,S��Bx9V�N%��)S��h4M���S��Ӄ��jy
Uf���Sټb��g�%�{Y#M�Pg}J	�@j�m�v��6�hx�7l����kҜ{�_����\`7&=����/UR����y(��^��P�!�[ۂH3>�C������� |.�B%~sT��%
�A��#��6�_7���XP�U	�jd(��3�T��P�ZF�R�Byޜ���}J�$B���]��H]�;���F@��!6=p�ή� �׉�b���#"9����w1B@m��5ٿ�o�t�Xi=><C3�*���o`g���NY��ٗr2��֋B��Ϩ4+��Wim����Y�����H<W��{�4v�E�]G�26%���/l�A�NF��n��M�N��H�1�̞�#�oc*�c��ϔ�5Afe��]t?�o�K-JV��$LKTp�Sx��ʐ��ߝ�c$��ؾN41�/����Hg �7���I�T8�#������a�o��p�T�ZjM��sB(��[W��_��4ⓩ`��ۋ.�����?�T��y�O��`�j�U��(�lW�B><\)D�`Q�Jt4c0��m�N��j�:	N�Da�@7�L��	8G�褂�x�I�1Â�H[�"�B��e̴����0��)�ur8Q����j�»"�����w+�"x���.&���Е�i��*6���ޝ`��U`��#���{��C`�r�3q,�'a/oZ�K�t�ovHŴV!���t�nÜ�K5�ʹ�.jY�ﳤ:��ғnr���'�����2X�n�X�!L��"B0]�Q����.�Ͳ:dc�X��:F�&M�*��b�"���v̦�����ܢh�����2j��B�k1�ص���d�0�նh��$����؟p����r����BS�}N2�[�;P/�J9妄p�}I�z��v�\��@�q �!2lv�Gm_/[�H��G��n��uUe���"闁����%�ۆ&Zʌb��f?�R���m������3i����Ca�Ǖ�yZ���y�D���$�o�Q����ܒ��e8�k<z@(z����i���MV��`���ä�
:ޥE�rjA�؃����.e��"?�0q������-� AOz.�֫S��6!.������y[N�M�ֵ��(M�X,AMy�J�G&��I\�C6���-�!\��ey���)E6:.�6	��{T��Ǯp^���s~�5�g|�u����|M�_�Q�����/J��!�!�^�@H#Ck�ޅr!}H�������S��:�_dJ�vK�b�����I#��}�/���V����������X��w��S$���v�.��y��X��ͼ�3RF:����1n��j浻ͪ�Q�|�y~m�;3�
i�Pc?<蓆�~�C�?d��ԁ���\9��u֓��#�\z�U,̅1�x��{x���B{�\n��G���������E�SW���q:�'�~5�}E���E1d�/�K���,��Hsoh�P����h�7���8kyH���R�6����G�<����^=���եw�tg`[ƻ�̈F��
��<���H6,Ӈ��L�PL��
g��Eɯ�)E�����}g�V�rj�8}.*3�����F6��K�y� (�l��1�=;�M$i4{A�2R���W��DWcJ͂������5��E��ac�A��/Ml�Pqvݶ�bz���@C_
k��8�v/���#�O�5�~�0��{����� %�LI椞Z��c��� �f>:�5a�t�.m����6�'%���r�RӸ��;qsRG��M �(��0��e|��&����,�W&�k�*a,��t,��������� ���\ٳ��T'���`\�&$�k(XR#�I�ߣ�8��g^ s��ԃ�����3o�Л�M���D�)+͛4�Ю����;�K{�@�3��%IU@��9�;��Q�.�yVl�S������� ��g	�R��쮕��-&�9���'��c�H�7�Q�`�f���?�k{.:�g������̨�	�'���[�?�*=	�E�}����Y��	�q�'��=�f��+VL�*�@�)Ią�t�%,��-�x1�9'��E���dZ�{�A���a���V��l��$��}* J��p����5���a:U
�*�M��d�E+�N�&�U�c���0!@:����.�_[�VDa# �J��＞:+�6��,R���� ��j'i����G��h����җђ��M�o�e�TT��-����#|SM��C#�c%i��Rܵ�wKs�"?���Aʏئ�G�'�'(�~:L3�@S	.%*�}����Z��S�yzI��a>�!�(�i�t���E�K�c�&QC$Pm�M;p��m".��j'���@���Ӱ��HZ*Y\e2ӷ�0*K�'h�����Br$1QgR���G[��25��ə����������I�:JC
��Y�|�v�B�W��s�ߞn�D��Ӡ�J��&.!�]��M��NџQ��N��ZI�WM̮y;���>��1�"8�9Қ��Ш?J��h���L�>2v�$�ݪ����Yа�{V���1ztI�z�Cnx�p����/M&�됙�3w��m*B*-���/Fvӭ�A6Wg�1��ۧ�xa��Q0���x�����2�V�'��2��Bħ7������� ��m���߰�&��<*d٣�A���w�3�o);����h�\���d�M���nAn�����c��D��M�M����#Ώٻ�X?ZzM� ��N����pk�?�Ρ�z�<��J��'�R#�i?��}�B���e����IZ������`�׀S��fiV1�~�� �>���ۯł(���.L���K0�=��_����I�G��\�D���C��[�E�B�*%���<�P骷��\8���(r����+�֐-H��8� @�գ��D��8�P�$:c�oSuV`q�L��f��O���S����*��h7�IK����X�,戲*�I�Up�r��
�H�q�6����^�wdM�űhy^!W�B��U27a��&Ϟ��}�= ���[�S�?���?F��|r��m����H�.�����Sf����sz���;���n���,�|����������h�ͻ���p���s�n�~��#�fﯘ�IN΃�y>ίv��#>�сݻHwX�4�_8�O���=D�n%Q�7��s}�W<@�~����|��������k�A���֞����4��,Vf��z{nߍ���3?�%���(��O�ԫ8����e�W�C�U{��G�M獞H�-�X�6���o�}x[J'<ڽ_g���A��$��6B��&}� .C"8��j�_Of:/�8l��;��hE��cwuYL[l���٤6?v����LWD7F��dn�{���_���D����xb���L����*Z������%���H�X
�L���+Pa1�0�V��+��,E��^�c��Fz"�ŨZ�gDj�!vu3 7�nЩ"�E��sN��-�;�듼^B�ګF��p*7�F�I˥^A�5�����!1�R�4�FC�rؒVZ1@�x��i�k�ʴĽ~v,�|yU��Lm5ã怩��7�է��dm!ŧ��Oy�8�t7�`�a<����r��ˆ 5� �aί<�ooGSH��<�L��������m����G��+GOo>�kP����P͏�z�������O�dřC@�Ӕ��4X�䳔�#-�I�o^�nG2{��#�8�7HZU��Xy�|��<�D�8 ��*e�_Ƶ���W(���Er�����d�UDM�7�I��~��j�y����*�-���Ѩ�R��9
A<�Q0W\�>��#���f����u��a76|([��(QX�)��Gލ/�%�B���-ݼpp�V�U���7����m���ȴ�J�8����}��~/l��@�6�1!��̰�i�$��F�F[J�+���,"T"TLNM��F���/�ί�:�+ZEN%X1x�P���-M��R��(f��NZ��/)�W����[k�0�����W�ʪaen�:����W�$���B���VtS��E��㵴y�u!�������飫�o1�fZiۺ^[O�S�o�z1x4���5�R�on['�5X�;A*�����R��6�	�J<K/a�=�f��*
����ټ�_��H�{��Q�ڷ�E����j�`���!��]0h8�,`��/�G����'�j�Y�4�	p����Z��(Tȏ/-<"w ��Y-�M���\����-b�]�q�k����J�ڑ)j�I�F�$A� ����ƃ�}�j�~H]8ؘ���.-M��u��`g�Ŧ�d���('3�x���}���"_�O_�j�RT+a�"1A�����ߦ��]��\�l����"�M�f&�@N�b�i��3��Q��5"��	|�,B���F̯�����i�yQ�G�~C��q�nD^#8�D����w�>kW�g oo>�,C�D����q�kY5���d΢��x��(`}�+Q_�9�?	ü��>F�9w��hB뉩��t��T�
��}����s�&|�w+�x;$����Н�[ia�R��t]s�7xVnP/��z�a3,�x$E���ɮ�-:U6�뻯�E�.�*F�����]rB��/y�Ĕh��{GWP�Evl�P��~L���Q��F�����XW��U{P�:�hZB�[1�>M�|aE�D��R^�@�y��XȈ����2�g�A���a2����Vm�*56���`;�菰3��F6֥�O.kE��m��jr�4��� �M%��-����4��͞�<�����4��ʐ=���'�o#1,'c�iZ�,���-�o�������a������#��<���6�4h��7�Wy��y<=�5}Lt��6��r�x���֐�zA��`�cv�K��������Zt(k��HU;��;0��p���
S�"��8p_�� ���˸�:~�,&�]ǣ���p3RZl
�k�� \�ka\e_�."�ݶ׍\�!*BѨn�/]��1o�+"Vy!���>ҝ��#���2����^wzOcH1,9��~a�巂��Je@
�<����#��à2�0�����4���ω��z#R�;d� |�_,ݹ.!��Ϊ�4â�q��S}�pGp*O+Kt+ts~ۂşx��������Ŗ:.�b;F�8�������7���qâ���eǌ�7�=Ҩ0[��˵��Z0l�w��Y�ܨX�"��	L�K�����1rTb�:us�"nG��5AD+~���e���X�&޷��,�h�-u]���3vJ*� ��{JwI	��BE ��`�#���(��.ͯ�]�?�/'+��
�wE���g����|�_1c�J�j�RVo�����=2���2��M�kGѶ��rkc0��itNl6�$��y�0�n����totZ�M��� ���M��V����U�M��n����sq�^�% �2U��v&���S�,^��=��mK���=������#7�\�,��� ��/ 	WAd��}8%�>`�D�)�ɶHΌ�t�?"Dgly�K=Uy{6�iњs)��\��ВkV���V}��ŸSY���ҹ��]2���%LQ&75���#33��0��B�ʄ��[.��T�=^�Om�>���
��O>�%av��O=���������lu��"`�\
����/�Jۇy)(AS	�)ޛ:i):	�_�<(��\8`{\ǃ	��O��c��^���~�C�:�,tx�����X����Fo6�� o_��������*�3��?�!]3�kF̅���P�hV� ޣ�A���Q�U�)���vR�lF�2&����	V͊�Ź�3��r��]���E��m#�Vlj��Y�ɽ�B�վh��ާX�������a~��q� �/�y�>��@�yIZ=C*��С���|��6���@4������󡍁<�b
���8iQK���(?�R0~��,��M�
�D֚�a��h,Ux�m�6�����Y�	�N��ݐ�d!�e�z��Fz
P�MB�[MD���)�Ӝ�:�SLҜ{$��^:J��E
s88�����0���FiqQ�֙��>��HS(a�N'��� ��W;��R�]�$#g�����Hz������k3��ԜN&��7���Y2����#џL!>q�/dx�P'=c��ɞǍE�R#:hA�1#L�L��L*$����x�8�迯�#J�<��l[�i	��4�0n,`�ey���O=�Ʋ).���[)��R��΄� ⾖��ptCMZ��ւ�����,�W}���3|������c9}��cClű��l:p�ݍ��P�4��@�R8��9�if��>���z%m�x[3i��$����>x�c�l ����0�Pn���+�=�ho�i�)Hw�:��.k����m��uB�f����ޭz��V�!|Щ�]�/<�d�<��t�ˎr?��d��Z����%��X�������q�h�=��B�`�����M����uW�S:w����1�u4�R9`�P�$�B�l��Q��^z�2���/��hZ��b�sX��}��v�����,����vx��%�Z�Z�M�~��ey�w�Z'H�9<Eʵ�@�nj�b���>��	琱��.Tnw*V,��ͧh���p���x�n�p� Z�����1��uzZ���>(o�;�5k��4Q�d�hN���c���G�,���q���_��@O�\t���$���f4]ʯx���[q�e�K���p0�̈́X����+c.3=l3�����pX77X`|�;�;Y���6�3�i[C���4Hr��ˉk&�7ύ���`՞���"B3��[��g�t�a���V��sf=�
����gZ:�ׄYh��Y �c[��99LE|�Ŗ�Aܥ���e�2w܏ ���������"�oK!X-8@zo�?�0�ψ�ӻ��>P�9�-H&�i4aV��A~ܣԚ�u��-�p�	`W4�ۊ�7gޞE�/!N����~�Y����_��ޑX��Jtz�����)��c���y�-�H�Ӂ㎕���L��-���ߍ֫�|~W�G����(���9�N[�/uZ���a�¿�d�s9�A�Fiq�>P���b�c�ϜX����KS���-�gsju�{�i���%�u�L�m� �S�(mD�W2�~vx���l|{��1�n�'�\�In����Ԟ��%qX�*����y�}_�t�[����P�DT�xÆ���C�F����G��ގ��'X>��X_f_�Q/�d�prlo��_�^m����Q߻�,��� ��)X�`��h�X����a O�������S�N�VH��%��,�
��O�eȕ�xq2�E�����#k��ջ.n�Y�K��y�o����K�s������ZioV߲�rd�x�������Х+2��r���_f�a6ՀFȘ��g�7����Hj �`n|�����+��[ک�R>1�Jc�1�nJ��o�m�/;c}?���ŧQ؊�B��������a�߾P*v��2~�q�H|�v���}*���}	{R���!�9@&���5 n7a�W��7�k�� �pW��
�xf�QB�jϿ��$D���_�ޘ�i-��q�4��}P>���^�@�A	F$<f��!<6��OY�(K�
�vf�v@�����܂-��o�,��!U��j5�a�N6_(��P�1Lٷl]�?�HG=� {Z�h��e�
O�N*�Ԛ�.}�y\?E�2�oRN�5��D�Mp"� 붢��z3p�9�|�ݸ1���C_�|u�mC���Ǜ���ܟ��Z0�a��SvH�6�Z��6M4�r��!\F�t�"r���clp����{rs�i�"틂�lKb6��/7&��#t�e�[��|#��O�G���Cց���T�tf@�P�M��kH�؝�KI:8}L�^ѱ��`I��!��2F�1����/v	�{$m�h�䚉b��1�P�1<B}{�vK�HhـUN������REM~���w�}1�Ȁ���ǗgcP��jU쀐�?�E.�yNؚ�V��X57���m:�����}{t���^�9'���k��$*{����;b��)u���ۭL��v��3"H�:k���\�+g�>�4�R�6��"�X@�03Ihk�7it�1�5"o2��-���W�߇�s�e|��L�O>���zY�U��7Yt����"6�J�ef���t �9�}̤�^.^#;�]���W���H�_��`�����c؞U
yy^�(,Y&IޮSV���L�@P�j��V��&K�Ga.���v��Ƽ�QG��8��
����z��ޔ�5#���𬬏nZ��/�s��
6���K�
m^B1�]��u�g=j(��^��O����t�6�c^���9R��W�ʽ��M(��C�AI_ϳ��?
C���̊��/�n~.:W�Qw��CZY�y/��ZƁZ��N�E.����}޷k`ͧB���hm�?���[��_��5$Q5S��(y"�'�� E0h����k�:�\P���#���B��bRu��9��'�b�9�(�k����+��C�q��r�B���.2 i���"4����?ۧ@m s���(�ӿ�h�Ks�&��E����d���T]�ס��h��f�1]�`v�e�[,~�+>�Y�nrMxRC/�i����;D���^%p�u^
s>��8���)�N?�^)��%?��&���s1��7c�$����v��vy�,r9�Ze�n�!��s�|�X�h���>T(�V�p[��|X���g������՝]s�S��l����k�	NV�k�@�X�?��+��/����uDN�������l�sx����qt��_&�+P�x���D���:QZt�sS������a������kO�܅�.�ba:��G��b��B��D.���>P��p�**7�)���_{�ś�yLxp���my�ay�a5x�]gh��
@� lj����L<N}�eV~e��ش��ǛFK�'�?�֢��"���jp{�Ȑ� �u�x̚"�_C�%�=�!�)���Æk�Z�2B����7��'�A�?F*���Ue��٧�̀lp'��J�-�o�������h4�k�S�#�v��*<M;��g58P燿RS?(�N�"�����>O���!�0���԰����vG�;�E�0��������� ��7WawV���w�ϰr�u�| ��&|�����Õ�,����V�+Pir)l��������j��4h~�!��k�6N�@�b���3��삺�"�{�4}��nfP��ĺI	���)B�Y&������z/���R���.�f��Z,?)nXJx�3���^�R�_d�:I�O�e�"��4wj�P���m�ͷ6ŷ�_�U�h6���,���z�K�s΃���]$�TKs��|q�Κp��P�f*_�s�k�V�`��ρ��DY<�]oF|H�� �}:�k���>'���up�K�Tڙ�4��7��$F�L�ڷ������ N�h�	��[���RHפq4�X�|^1 ��N�	�¢�j���ym�hE�e�'����&�H��A��Td6>ϿQ�В��!zL����l������Տ�i�/�V�;[�A��� ����>C�Ӎ_�ë(i�ݑE����"�#N|�>��?��c��>����D�a�Zd����Kt�H������+�Y�ѣ+e��o�S�n��o�.�&�1d���5��{T0�
l!žqb��f��d��-ۅ�����`k��1O�%�D;~s���a���!�B�#������:1v����4/�pޱ���7��	���~3Ĭ����R�v����#��0H�=�;����T=wT���:.�b?�4!~�"o�#�l���4���fM]�e6�G�g-csK*5Ӷ�Ry����<�}�M����h������2P�lK:���Ѯ����zUPI����)j?�>���+��r�յ��Jq���9@F=~,.ro�z���%����_y4/���#e~����ێ���Z
��Gf����r1������s��u̇�W/��'nJ��|$�mN�n֍<7��dZX<��<)���������c�$xq�Sú��b��A�`���*u�V�<��!��\[*O��d,���y7�V��J��uj�"�D�>y�i"7�E�"�H�)�4(������O}D�zפWb�=Yߩ�j��l?k��Q6���n�@��0/A��z���t���l����ZER�J����NIfѦ���]�l��m�׌�m�4;�_��G�?ނf(`���1�:� ���zp�r����}2��?���k��m�t�&��ϼf�� 8\����ԭ�7OlUm��^I��B��1����I�����2��)Z7U&�.�F`����k "�B q׈z�1��4�O�k��(r�^��1������O(�Ge{2�姡�	�v��5ͫ$�3�<�q=]����-�:��aG՟Jp�|r&P�ܱ7��� q~#	��$���&.�O�g��:Ӎ��B���T	�N'�q �C"�@�Q7{l����b�����o����@+' p�g��I-�����F0w ���ڻ�F�keX!y�q���p��>�hqt��WgW��<��9ע�2���G�Y����	���4$*�/����܄��)R�G���>;�k/�5�	�+�?�	_(���j,Zg�2���Q�Xּy�w?��բ 9&Q-\B�o�*��¡`[�筤�#\�P�Q���5i#�����ubc�����6��3g�:Z�$����l��հ��q�e� ��
�N�ڌ���ʠaj����U���p�,
6���y��iK�A��v�(N+#3�LU����F,!��6�r�a�C )7�<=q�5�� ����{Gp���AnQD�������k���n���s��}���U��h��a�x6t�t]/_��Գ)dd��f��RW21p��.7�NTf ��,��4�ݬ������h���u���O��1pq�Ѿ҄���j����H� �5� �ډM�����oK�B���(�i�v~g����
��a٢t������&=��{:�b�t�Y�)l�������ތj�����a���cnЙ�s�}:I��H�5{��1KG0�W7��f�"'fu>a폷& R�mn��~u�7F[4,Pմ� }$��t�%@��o�{S���M[,N�z3/_	YHM��>\j�q�W	V�@�"#?u��Y�����г��er�9�ץF������l y]ۭ}�騍��WJ3+8��{�vx6���Hz�D��:p��q`rzx�64Y���"v4�Ŋ¼�"�a|��,��qġh��z
����\����Q�꿝^ma�ME�.`����f��:_Gc�Ē�U�J
uݸ���~;-�܉a�+��_m�Wq,ZNN��FFx �S�ĉ�Ԣ�v�.+f}Lu��7�ҧ禊�UQ�xL�ԆZ����<�Z�&y�,|�yXmLʝ��=�	%k����!%�'����dtu���m�_I�[�����U�sL��O{w"$Ix����/��z�T&r6)�L� y&E�j�> �aB	��w�J=�`'��0F�g	SF������c� ޵���S*��t�\�E��y�@����X^*��P�vJIS�f��ޯ�d�R�6��실	�vs}���o[w��|��p/����u�tXψ�8%�Ӫ�U"�ND<��	|�a ����*eR����������O��2�%6��ߊ�g�I�x�H����s2����B���rRK{�OB:�v
�?N���}��R,��E��F��g��듰�2oe�2��-Ǭ�`ܖ�U�֛�X�荑d ��^��9�V��Q� �\��6��:w�W�>�G&<MH���9��L�(AM��>��0���] 흄�ֿ��9�`���.L#��ƒ�:�g5�����}R֗n&>�G��LuV��&���]�里�;�q�Y�azr��]¹��9��M&��$`\�:���L��c�J��/��E.8 �p�;���/v����'�{h�P�]4��:6}�;���B�>Β2@�S,�qEؼ*mcx��#�1TqbäP�Mi��ɟ��;����l��`4�yW�hO���9g{�{��ޓ�d���L:�o�������n�$U�"Uq|��� )ߦQ����5s�����U��*J�6�~��B��Je�0~<���"�w��b��AI/?u�
��㺧���?2��~�ha_s(�6�	�X�[7!��<�J�a��z�cf�(��^����_Ώ!��?�FFAqg�6�ֲ����`ϗ��ma�Eէ\���v���t�*|�����>��(DTM�s�P����P���'f,o(k2>�RxZu�ڤ  g��>�������;&&�|�c����1�)1�I�����Z*#w̅�eR��LTe"��XOO�{�*#4X�9����=p����3���ا��\ ]���c	:�m��=�~�&����@�@êq�+�H��5��g�����}S�74�.��5���bCq�[s	s},е�4ԃ��p����7�y�Z�}�u�>�㞧~��L%���!=1�CL@�(hM�ؙ�\G���ƍX�J�k�i8�ǎ�e��q��|�H��׿���9�G=�#(�����m�;��_�<	��5�;��<At�{�mq�9�;�z��\�k�j��=���-�b�v@n�5i���FN{bu�B���VlZo��=����!��\2����sf��a��xu� �(��*K- �-}��1�v'퇐�Q��@���'��3"�8���;\[lO�7I�&�����g�Y��(��G��%�2�;�}�I%��� }:Ly���s�q�)���ѲC�5b�֒��j�>����<�v ��Z������؅iߑ�̀c�_������K�;/8�?I���n�Xv���$��K.(��2�}�MVk��_.�lT��[0v���(7���adh����{֖�r:�cV����}"����1b~y�ƹ��ࣈXXΫk�ഒKgÄI /�/5K%���t5c��׺��>6�8t}Y.��.S�&>j���_�<���>��m�Pfe�@U��)sU<�z�z����3[K۲�:!-zy���J
E��7΄.Y�m���I�ۓ��gѤu{�mD]�	2��9�:ͿUl$�t�b����KB�:@ܠ}�/�������\QX2B�5��뉠8mƆɱ'�̑nQ����_����G�m�-����A;�@J�I�gU�Q�'�>�w`�f�����X(��&a���\[K4�z��-i�15vhO�9�
'�~B��+b�?������y1�9�A4p��oR��|�kj�0Öi���u����K:B~n��T)̳�u��P�N}ǿG���2-o��3�����[�A:��z�+>��WҀOE|�8�ڵ���fE���Al�n �8��:���k���O��:IJ�}�r�fCF+��V��(H%���h1���rX�V`�+��"'��9�@��6��)#��y M�s����ֽ�=��WC�)�㹝$-T�.π�!���'LKWK4��ࢪ�����%�YQ�	۩妔
�{5]q ����yi�e\���oӌXN�m�ïe�C���`mi�E��?�XΙ]	M���4�)��m�#M����v3Y�|����N�8ͦ
��v�^�R�a�����1�E��(�w&́��
�qZ[3C���P}2�c�6n����t�3M6����Β�&断k�2ZQy����x��i*ڤ��++�J�C��/K&+J�\�-G���IT��n�+�Oӱqwc+l<׮uHb�?�|��v�0�<S������5�8��'���� wD����=5������{�L3U�Kț�ږ�� d�ָsb��1vʚW'IR�(��Ά�$FI�!;��5����׎D&���K�v�vs��r?�/ ��s��(}�Ro�w���)1�#�u�y,������<s���DmnQ������8D��{�g0~h�	TN�?��:X����C�j_N�,п���=e�T���6�y�Kg_I���{LYJ��ِ��@$�C��I���.��3a���������zU�(,>�U�����9P������w�lovP�9D�<�ɒ�)yU޶�1���~��5ov���8Io���c���>d�G�MOl���K� �v3�I���O���R�v�,捲n.]Y#�O!\	���'�u|Ni��7��gYf�y�����^�|@!F$�䶸��M0��&���LO�Ff�i�r���/hrɂ%ת�a��L`�������Ŷ�GD��P��(&�9[
����om����>~=���u���i��%��N y8�i�s����B/W���jOÝ�]�21aw���N�VZ�V]P����2tjo/���qĂ�z���3wXr������
c:��h2��Z.>cP�H��3e���@�\�R
��2w�	�$�?���F}Uߦ�|V�s܃�7� k��\Cj��p��U���u�9�����}% ��@��>k!��Zu2���v0�R�RC� F[w3�n��7��an�%��p(�zw� �����BEΈ���a�#f��ڥ��f"��v銮�N�_o����EB�o�,��'E���4�]�%���kiYC`Ͱ���
"Imo��[��Oz���ep���	�oX�L3�q�!������Rx�C�#��2��+B~�z����rG�W���y��j'��j�������S8aӏgO�+��5Z��\���Q=x�S��Xi̎���}`��oAPȵUZ����̞�bQГ��<4���\6/%��Q�r��u�j�P��h�����(nޜ*��sB"��^��K��h�|�8�	i�T���\u=\'V�̣'�1�����?�T>z�YG��T�W�o��u��Z3`���}��~�4�d�qڜ(@��%f��C�%w�|��oM�7�y�Q�p^�ul��!���}/ߢ��Ca�=�����?�J��FR�4�,�����dW��zˢ�c}�9�6�:.,���ǗW�)�N����6&�F����p� ~=Q�Z\]�ӟ,����7��O������,ߵ"׷@l*v�6!V��/&��?I�M��m���d�[��j�Z)>�i�˶�E�ղ1/����Q��q�ӛ4�xWٗ� �r�=��/��qD����c|��.9S�D��}|"����QFF��c�����ΨiS�J�\��*#��i� B\����K����T�q�P���:)3���D6"��6�F���۶���p������_����[�[4J¢�|�I��B��q��� L f���V5�f���θ"=�v��OgpTN�r� �L�*��WX�����X���N�q@XI����o�^U���V\ߵɔ�@�GVj�n���%��-��ȹ�w��-�^�� $�,��n�p���G����3�뀼�E�l=p�,~�$	8�Q� �&э�_������3y޿��7�����	���z���]0CG���ѡ�>�tp_]�02q>2��:sX�c 1��'Au	��u:I3�XX��(���#0��lK����f1���-�c�;K���,�Qwϴ�̓g/*�r���������K�5`t��[��~Yzve���s��t�}5��B`����lc�����)`������gr���M��^�˼�q��r�V�H" ��޻�8�/`C e:+nڻ: M�7�0*6��zB�*m�#����}i�-(w�������&��O����G�E�W��`��[����m?�'j9տ����@�;u1n3�:V(p5_�"��{[���	`���~c��B�1*P��V@��ཉL��f�7IK,"^Wh�.{�t��B�!N�E=���P�;MHXw�Ίfq��ѯ�r'iK�ʃ���^|���N�����߭�Hu�/���Q]��U\)�?d*�g�e>U\Q(�z
F��Ƙ�����)���i~�n��B�M�RT�@г�M��
���:��w�>���yέ�� ��A�W�D"9�0��GN�ڏw�e4*_	 33=}qJo�Ӈ�-���W�����渌rǮ��8��Ӌ�mޙ�qEǅ��T���ЖyK��3�D=QXQ�@�i��G~p�i�7�/�Q��xa�jH�{��U���},}��;Ix�����rCb�|P�$�&���B�aNH��+c�6�x��囀����_�v�!azWj��X�3����*jӲ�^��M�x��ޣN{���"�*������y���
���i�2Hҟ�\�7Cͱ�`EyP+>b���������bkʰ����v��x�q%�[6|�Ak�� a��⺗:0`J�+����M'��TV��*y�W�7�" ���[�{#G�DV��l�����'NW�f#�;�(�إ4!��h�"�q��}�cb['�0��J�M�8�t�������}�~_К�뾿>�[�i �%)	jY���xj�F��4��o^p"�n>P��v�u����7���gSj�G�d�.D9R6�%��d?�֌N�Td6ҽue6�6�10�ع��B:���y�+�q����c����篚$^x����fm��i�>n�G�㨅
S�;�(WS&�R��OC��+�`(�nnT���|�/������ϣ�,���}��1����s,]�)�'ۉ�~uJF��2lӧc$��|��kM�f����Y���F����<�l����quJ�6����n���2����T�9���b���z�Co�O�^��G�iv�����'aNõܔ
/�
��L���Q. �8Ѣ����k�u��\�&dO�{{�l��R(�Y�M�������ݪZ��,؈�1����)���2w^Ґ�Z�'w���َ8���0GbV2{S�����1���Q�!ħ�=��_�jE�H��V�A ��~N��xp1"U����Ub9��4η$�B���f���Z�tG�q.�۶_s�{^��$�Չ�krb>��)�lX��/�'��@�(:�my0�)���f ގ¿��Ght!3�gʮ9d��iĉW�R�v\]q>�;9k�Z[HGD�1�e2���Z$��o�my�SU�-m�2t;��@#���Qa��}�픫(r	�~����� ���NEdm/j~"�)S^�w����/��ߛ�4��p�^���5�q����I��}dt��9Z9
L�(䞤��u��bnd�N5Җ9N�"'E{�U��w�Ҍ�`�.2[�7��n\&�[Z5�H��U��{#e�y����ӥ�Sl:��8E��Q͘�E�p��8��z�����:NbI|�,�\�}�S��h�G	I%!hfj� .{4m+_O|Bu�Q5�� "�� �0Z�"�͘�77^�aW������!�Ef;�֣����_�����F�g	���w��9�|�)}�p��!�ٛ��?��i��;%���\x�5F/o���ۯ�R�\q�}vj�p��q�'�͂���z������,K��
����_{as����z�>�GfN}�	�i&�u7$ ��L���f��*�U�/��a��4�w��r��u���u����`��UJ�C0�>JAm��復��@hp�{DoG�l�����v:r5�e����+����Ie��0��ͳP{s'�b;~�D�to8���HOn&�˵�a�q,�0ۛ������=���
���(u�C��8#L��M�w����B�ʻ��:��
٠1�o{��u�&R�d�\�A�@��(_j%�>�%��y���9R��nlL��j#�|�۰=����͙?|>nވ�{{��1W��r����j�P�ȗ쭐��ᡇHr!��ĻO��V-Y��������U��|b�=�$MW�ɽ�G�:��<��&��5���q���3�;� ħ���T¸{ly`n����-B�s�r���ޞ�zG$�Wv����×���ZtS�V֚!4r������[���A��n�qs���cס]RpFV%�W�я��f[��D��"�P����w��"v����m��]Ha�#�@%p�{�״��d����T�D�9y�T��	�@�-�Pܚ�����b��d��21-�L���Jfn%0n�y����-�A���[�:�{+b����w���#����͝9�F�K�y�򜼵��AA�o��e
��Cc�Wr5����;+}��A�?�
H�v9Q<:?�
�-�C�0�oo	f��;5o�DQ��@�3X���ɛV�8���n.j����h�~g���#�"6oOએej%4)|tc�M5N)7=A^����h��ci�j;R�f�i��s�mq��*)��%JzvI�D�> �ę���T��/U��Y��U콛�������MT����摽@ ��)���y�kG��D�l+�) ��(���F�mT�ŉ�����Ɛ#�������{E �k=��{W9��H�a�P.����~����Q8%�u�i&�H!Q )���M��U}�U��g`���4͂�o� ��������z JT4w[��|��=�ǉb�h!j���+,@m�#�D'���̸geG�_h�g��>f@�� ��U���|���m�=��ˇĜn�R�F�j��!k�d�N��3����p�5�S@%�
�d��a�
?$#��(��6�V�΃l��3l�$�'.z���ɹ���/�&�dH��2��eK2�q���v������ �F�q9�������=R��>3�>+F����)��YF��AZ��x:6��2�Pos�s�y"qh�l�g��B���]~!v����z��ޟW��/�-���p�{h�(��A�d^il&,Vr
8	k�n���I�4u�!���w��ݒ�d���>QOD�I r�p��#�j����2�t[�Z"��q�)⍕�	�C���ft�y^?f���'Y��R� C�����ZOd�0�,�m6'��6�a4�t'�i4J`� �`>���Wq���!0�%�b:8�$��L���������`�_Ӟ��ʸЧ)5CL���%���Ӏ6� S��|��rˠ��W�MT�����摱-����=�'�>{�����������^-0!��:�S���I�K�`N4������P��X��N�.@��tJ����cF�q�;�l �?�����2�C��-OZL����H�*vm���&�,]3W2�0�<d �_`��y�Sy�F6�o�&��O1z]w|�v��1��ܐx���ʐ�������@��@���C�a��֍�W�-m��}d��9Df��~2�gNF���PzKF�a��T�T7"!����/��
jK�3�I"�kY��r��?��$��G��GT?�,2U�i;�QXw�G�1}<Ƒs��	���!bEJqZy�I�j�4�3��Dw��%�UI�
�'�_��2�<����=����<w�t�6�Q9�>�+��s�cn��y���7���������G�2U-�c��c���v�1��B�ڊ@]R�M*6WjM�U�SĒ~[��(qs(I�ھ�ZdE�e����v�R&�o,6��8)ڌ��x�>�S'�[��"�v����}�����G�8����V3*kz�c$$�����k��ʜ ���*Ǉ��nw{��r�}x͎_l�x��G��"����֡Î(J�m��fV��58NQ�ӌfS��m��0Q���;N��Ȭ.bZ#�:�2*P ��D�as�,���f�L�,���}�	+8m�w���՗������%��粥���1������%��)wF����sc���P0t@����j��%5m���H&G����w���q��j��b~ =�����)-����̲���gs��ۅ6���s۸�/j��\���2!V>e
�S�$9����f`'�6�o��C�Xq�9`�4�?=E���f����/�����q�|zp�wjoj� `z��ѫϝ���0��A�s�`b���@d�M�h������te�_��z�~��Bѣ5�ME�L��A.� /N���{7'�':�]~�Mk2ؤh�Y	U�9�v��z�{(��q੃��)�d�@t���@ע
GB���l�4��'�HiŢ�ʪ����0��fA�k�	�@&|�.��4��m��Ĥ���V�I�z�&�h(S:r�e*�x��z��#�I��°OV�_� ���h��ղ�-_�����-#G?] ��5.��[@��JѦ5a@��s�����v�Q+%��:�,)�V1�\������W���~��)��8����[���qp�n�k8���<R��6[닅�����V���l6BҲ�tFK��"��G���8����������=K���������w��x�82�)î�I�&"r(���b��9b�yG 'q��+d�#B�}� ����EUd+U�ֆv���#��?A�gjU�]��5���4�Q� ���]k��/F�L~���izL&$-u�!��6D;�G;�B��v ��@�.�ŜA��ek,�5S��H���2o1\7�*���!�������y�D��EW�c��l<x �)I�83�3Vڙ���y{_� �3"�i	�Y~j�MCQ��k�2G��y@���]��?�Oa��w"��d�wt�d�\2���� Y@������HɎT�$���(:���Ab-��i���)k�i��P�S��Gp���"ҍ� a���̎*�4�1"���^n��3z��R����4���Rᵆ��hZ���Pqã��#�aѲ��38�֠|�J���=��d##�Q��|tT�!��5+�x=���Όjyk!��<�ɹ���Z��/��w��V	�̊Hh�W�ZV$y�Ć�,UNH�uH]�B�u���t���,����+G���=w�R)5<�Z����zs�If1�*�H����޻��]�x��2�w9��-��5�o�������Jy����_�d2xK�!Z�o��fE75����k��<ᢍ�os0�/�O�?��܆�B7I��&�B�����TN;�e�-�G04хW7�+3���my��*���>8����o]^�� k�㬬2��Sٸ��2W00��顷T�5�o��a����7�Ҕ	,|^���g�(A�� J�#�lcB�"������W'�&����x�}���l�Ns@�n�(�U��&hAP>= J&�W�Ѣ��똇ӴZ� k�4���㔾n�b���93��NmK�g!d��O6gP���N���6��YkXP��J���8�	�SO�����3zFyC�{s[���3�;x�˸3k.�;�CS���S	��T��s-�0`6��s�	=���IhV��l�-)I�%�@�K��L�|9,j�Ih|��`K�Ckϳ㾖����F8��_��Ё����T{�}ӄ���L�����֙Ȗ�� pm����+��hv-D4�ٮ.Ԁ b��>�v��L4aOp�]p?�6�H^l���0,<��!U�஍̌:�%#0�x��a�,7��l5F��瓾Dn�V�NIې E�Gm�(�\/"c�c�Y�D�B=IH�Z�^S����_��Dp!�M�M��]�Ja��{zF�5�z�����y���?�~O�ޔԛ��ڮ���+_�mM�u���꒮�0�g�t�G��Ť\?V0 �Mָ��,�%��U��SȘ����/���r�f$pX/��C�MK��h7��ؗ����@(�����6�S�3"EBfu�b	��Kc_zz4��?}Q#���!֦:���=�𕃘�n���/���4{]��>�C�waX�w<�_��,) E֫x�)�B.�b,�d��'e{��I4z�_I�]��J^E��
��%t��LX
��j{���[Q1@>sٯ�y�-R3�aJ����t$6$�8a�vBY.��3<6,0zbz��>�'��d�j3����f�7��m� �LSB�����ߤwaVC�Z҈����w#�{:ב?��kyBV̤�W(�E�#�B�Oh�i
>��L�n�˗g��o��_8E-�Տ��:#���8���Ǹq�$�m.jz(���-H��K�Ό��pZE��M�iv�5�È
=J���+��H5��Q$rzg���J1���Xw�-9�2�5�H>����UK�]7���Cy8��%�I��r�?./��gA��-�RA]).�.)2������Ѱ�|{��e��2OA�x��P��7Z�a�U}���z�UA��a2��:4�v{Q$��8��W�����3�̊s�YR��As4�o���f�=�_A����)��x�u�UC��r�^Y	uX���P��d捷�5�LIş�躕`��sfܗQ�9K!���#�x�`6:�.����Q�?��XWXc(�HiI�u6b^Nr!��}�;�r;�&��Pǚ�~�?��;�pգ���WvrL��f3-?ѪXsDm�5��{�<�W�[M���}��~Wn��m[}�|	��I��t=�*�I��C#Sn]$E�J�sm��1^��|sJ X��RA����U�s�v��l�(��%���p9/��r���a{l��~~4�\�����c3�P rhOՀ+�#u���H`�Z;!��o��*�ͼ*�j���.B�x���A�?���a�<j�v�@�G�۩��-�����<��Oo�����F��Z��#/��'ڥ	��?��;�Ey`<�ģ�|;y�`�~?�{�����!�o����ݔ�;֫4�BE"��K�����h�%�W�+�y��P�RV]&V~�6 Q��5�R�1Fb�3����~�-�N暳C'�@����^��Hkn����T|����9��	3RO\�ڕa��M��|�p�����5R%}���g�������R��~$�ҿn%'`w�s����k���*����i�}���_��3x� ��`"Ǳ�ic���{_w��P�֞㔹Jq�8Gn�!������7z�-��eJ���p>�Ġf�z���ҹ�]��D,fUK���o�D�#4P�V\����]��H"\��o6_H��j�W$�h�ht�j��:I������A��x�|�Bu�Z��Y���M''	hn<U���?8e����I�O)yA���\���v&��
ݗ��P��~XG[�-���tc��I���ۢXǑ"�{��SCTQ%՞���Pχ[�/����U���#�`&%��(av$����s	�]G��C��![yJH�/9 �B�f��݃�+]�p'�����Dw��*����|��S�!�� y�Cq�V�	�_��C2�c�|X�ee��L1`�����Pc������N�4���)���nr�C��OX�����^܉hpQF)׿0����:o�^GpMBU�~��}RwDR��vVL����fq-�B��OC�ʲ6��1s����G��~�xĳ�NK����٣���4���_����zm��1fD|��H	��)=Z��>n�/+
�^C�J���y�:�x����Ӏ��7۵3��$g��_��'@G��9����o&��Y���*����+B�{���0��S�/�=}y%g�8�}���v@J��G�
��A����g]�X��X<��Ӌ��b�O�PP&�XXv�C�f�a^�����0��A���\�-vҶWBSE�%�f����dE_>���뵟T�8�pS��D��;ް�����Pź�߲��P�qUc���?�"�gW�{����nL�H(�	�`�L��P��#��|���єƳ:�~��B�x4'l[N��^�X���t����+]��g�����tTI�����i!���U�@�MZ܀h��-rn����L�S.*Ύ~�ચ�x��F�q`:��p��U������wwY��!�Aޝ�v+&�Pl%�&nY_�O�_�*�ҾNB�
�|��q��O&�j�b����Co���	f^��ixð`����i��)K�W��R�o�?(a/{�����U��I߅pu4�D*&[�kZXb%�y����͟�[Qa�UPq/�ڠ�D����^����8O��:hʴ�y^?��m O��D�g�k�m���ч.���=C�^�pu�-
�uΘ���Y6'��o,{Ӏ~s����\ؤ���{��#��N�ƈ���7�V��>�����>��]�S�N�������-��M�$,q�kС\*wڵ�@.�ϐ�� ~���3 ���	������?	!#�A����[��;��T�O���-��̦�@������#Kd~5/�)�˅���\n� �.Xy����r��3�ToD�m�hf /�U�#s�A= )�Ƽ�C�q������W�ĸ�H��٫�d�Q�򳝯�Mcј��	�(A����L�KR��>o#��f�]d^o����zA�P�x�Ne�co�]3&@�D3����M
1�M�;5Oa����L[��֨a
ǉ5@j�Χ_����I�.)C&`��\��cu���:#si茋�S�	�Q?����	M�� �k�7P:
|�<<�b�]	���*W �<XY�x�<���`�ڹm�#G)s���Hǿ7N4�y��K6�AY��&�m�>ƞȬ����鑵r���X闔�GvaE�P!*UL���6C�Vo��^`���x��"�k�x#�4��i���MD��<c"�~�\'����.�SN�&�� ��r�)�E=fU^��r�V(9�������!���:���ё ����s�ոv��Z��N�Ӹ�gC�[!�8�mQV������khs�	�n�ECw����2	�<�5�� �1�����";B��K�m|������g�tm;����&�7(�P2	���8�ݯY��7Fڟ��K��-$E����_mN� ���)��ػep��)=��
���z��b�h�Ҥo�g]f����שW���J/�?fn�IÒ�W��Z$���Z5g�X&���h��i7E�h�{�۪��g��WBSsgp{5#jɨ�8]^/��Q��@,�������u�R<vW�ҙE�V�/��:B�l�<y/�1�O����#�'��#�45"�'u6�y8�,�\���ޭl'W��2떀�!(�<�j��>{�Ȫ�I�ɕ�#�ǈ�dq���p[��M���שo �`����dlgc(����3�����w���nh�Z�FzҐDvf60��;���N�1��0Z4�9D�7�0:��h���N"U��)�[89='7=��� �����G��ss�a��X�9���G����]�`6���!�ܸP��w�A�8�n���7P�8/����]�-Ϫ�i��ȗ�zS[1�na^H.Z*�Ee�c�%J�8V�-����N������s�8��'��Z�������
�ʘ߾M���`�����&��q����}dx����}�S�.P�
��Dq����}Hr&����h���bIC�ڶ�Jt>bne���mM0����ф�X�
�n�pTSG�ﭮ$���{�p��p[z4�5�âb���AM@KV�8��%���!���K`Q\�3�P�Z��"Jp�ac:�b�ٻ@�����!?4�� ���uP��O�h��� Ѩ�3��ߣ�����8g�-zP,xk��+���߆�~��O�Oc�Ԛ��M
���V�:JH��*��^.�[g�R{�����G2E��X���ѯ�%/�ߘQ�~|Ivm=y���E�NQp��}����Ds�Ցjg�)@�bhp�B	N,B��/���FV�h���[�{Jʿ�����9_�S!��Ĳ@��@bk�v��Y�ָX^����
�w���|���V���؍c����R4�bj:�ڲ�;��3i�:��f�)˷LQ!Xx B���*ēV}f�����}��k��^]e{���W.�G��0�F�J"o.�?q�r��)��FHϔ�ԗ1q��B��9�������IX��Qq��3p��0�@���Gd��$�G�^��UnD)|@S&2�o��ȼ��i�	�D���%EB��^
�J�m��k�t�R�����a��-�_�� ���N��Z���k9����ʵ�mqlO0�!{��hZZ=]ug-�+sh�?Gg�~�W'�&jQ9�hᥙg�tj�4�/�m�*P�ZDGt~�"e�>�A��|�&����[a��a7l��zk��rH�1/~���!���,d�<3FUܚ?֋�Js���[=�F�����n<���(�,�j�'��	O-qS�5��8�&�\F�q����(t��˄٤�����ҵ����*����9|:�!v�c(�q��(l�	���8���Ŗ��y*�|��/���7e�9�'mWƩA�Vl� �\�1ʄ��##@�������F��]�J��Q�Ӥ}�!>ǥo���k5~�7k�еv�pJ�U����o�+HF�0{��.�D*PO6H�v�\o�X�������P+�E���{�{�+�%��Bl�Tot�|�7��@����I�&j���TMWZ$-j	�����,��ۦ����H�b����W0��=HP���fS������3����_l�ύ���!����1���ɠD<����*��jڙ�R=�l����<b��
�IW)��%�X�$��x��β<\�ȫ���ǂ�U�uA�u�<��26U�QY�G6J�H�'4)���ַ�e7ل���`�V����V��\�2KЧ�>z鰲zr�E�6א Ku\z�?շ	�1��w��P}��M;�����v��IA�qH�P�����h�ꚴh���5�H	��M�C�WW�_�#�ԇv��n�5,��['�1�"�e�g&�a@��4����!/�=��OX��A+H?��õO|����.w�!(B�y5S��m�mx��1;���C�bx����l��N0�K��"鉹W���os U��60TwC��u��K]ِd|."�bػZ�:�(��| Y��>������]<�m�g�S3&<0x�!����}و�XA1���s�	�i�[�cQ:(.�\=v����A��r�x<q�)Q9���k��!� ]Pr�ǣ_���#�]/j)��9rb��q�6���C��\���Z�/C��
��zF�f�Af���L���N?( ��3*#�fMnZ��"�sR�n*�2�4� �-y�lu���!~�[rvEU�+��OZe��g��k�n�:�{�J�}�2���ܒ����spdW &BaVo�]�wM|��l���+`��<�~~���i��£Y=�/BO�����%�T��;l�㡶ꤖ�_��/�w�&��GV��E����b���7?�Ϣf�s�Mt<�Q�\��Y�R_n	J$U��;�gjl����=I$6��"�]f�_�%���z�>�C�d6H�U�!��}��u��&���}nAG���UͿ�@��A�dO�Q���k�{e�čȀ��!�xb�dX���H@P�m��'����+�i�!Ii]>�t�:�?45|:�g"�?�{JwDA��JVP�����J���(�ء/ټGL>���C&�g�m}m/��� �ʔvWCL	���";�F\�kǓ`!ë�$LS�@Q���N��\���h��s,��t�Rl��\%<㡖�wڄA�����FTr��Æ�-נ��C�L��}��6u0�Kz��G�F�%.�%Z@��#���]�N�L�����¯�lϛ���pih��&�
T��l��qHt�>���iH��R�FN�)9#�Y(��'�^���!9��.Mo��13>�=A1")���$������5��,�d�W���U�!�+@�W��8���Dƚ-K�<sO�x��!�+B�%����
���_�:57:p�s9��_��e$�Y��DU��>��D��gC�s ����WK�MU�ù���8��Z�6K`|�q���H�YmA��aÈ��Zih4�"��p���� C�V>ΎMB#�P�~f~��ZnhY�
���j}`����E}�l"�\�;�3O����Gmc��.�Y�10��n@���݆�������5Wu�രhz�b�/%�K'wQ[!a,^ڱ�ȇա#�O�����B��.Vh��gj��I��U1w�r���o���0��v�X�X脶~����\A��͎Z�k����ۤ.	'��tޖ�!�\�𥮃��B��S����#��H��'�U�-l�%w�W�+���:5�ˑ�|���
�g�j���	:%&��/� b�?w{]?�ǔ�I��^�[_@,,�$��*ܠM�x�F�QüJa��N6��ݧXkzu��UyY��@HY+���|�Z�TjAX�$�7��g)nGv�_D��k�X�~ty�����,9�o�Z!�-�1woK��}�j��uh��%Ԕ�^@cv�m���+Ф<��]�e(����i��S�T�,��R�
8Kuh�����((������l	�5�j�)�c`Qw�ӡ�R��<~	������F�plk��1���ç���Թw�x�@O ,V�cc5Nv'!B��n�DW��Y�r��kp5š��5�pqW� �1wÄ
 ��R~u�� C�����ek������ŝ��Q�Bg����p��`*�0�5�Dc  3m��j�Y�a5�B3�iBH4nK`{��:�ġ���̿�@;�ܗ�/{�PN�M9�%{p��+H����Y��K���> ��c�X�8�������F�_�u�/����a��f������ڛpŐZ<m�0#��i����ߗ��Z� �/����
���$�䐤�6)OQ�	�C�]�f��P��1�"	��0���a�t�%"�������4B�P�Q>�f��O/����D괱�����bɊ=�0�>����$�Y��lO��W�2��0(!۟�1�T��a����B�V��8��z][t�e��4�<\E8�[&m��,��;�L�W>��e���VD3�uK�����Fw)�W#��CB�/��]�b�s��dj���������~�!�y�M��-o=Y��5�
sY��*w��W��Oqx�v�R'��K���˓��qrI/ ��
+n&���w��M2@tY��I�����Ra>nԈ�L9��ɬ�u$��{l��֡���u���\�y��c�O76�y��#�P���U�����\:1*������Qe#vH�ޱ%R�)���a�³��loc�"L�o�r�^��Q�\B����}Ny�������Io/Q�����׋Xl����E�a�������,z�xI��
���������Z(^\��s�2�GU-�ٝ�f���YqƗVQdq�Bt�ԗ迤��ਚx���/��=���m���&0l�q����ԥ|4�Z���L����r��)���H9�g��/q�i-��ؼ�%N��u2η1 �BƬ42��E<���v����\����٦��aI�WP�i&��B�"�J{~��y{u3�h�O�ƦUay>��2@t���5,��K�B�����@A�u��h-u6�G��])��� �Gi�}J�Mk��A�WbY��3�;c��s.�(��%v[��A�f�Bh�� :|�M�;o��vm y zS�?)�64�1�/m"%�&#��	߭�lέp�Z��}RMt͹�!�m["v�guZb���iǖ4F�{�/��-��9������ȣ
%�m��j���v��:��e�Bx������Sϐ,%�{K���InjQk���b��Ŏ�0j�{�EQ��q���3�!�,9Y��r8I�`h�*����[6��'��@�qz�׏���G6D�%�׎����ۡ�ݫ�A=���+�_Z��-b$1dg��
�c5sj3�l�G4c���f^�u#�Q�C%���~iZ�b�,;
J�c�r�݌-����R����ic�:l�u��˱���k���:e�`�$Ǻ��XM�V�r��x'R/��������Zw�;jم x�M텑e��E�b�l�Y^zNV<2uI�Zꇗf�|kb�SƌZI띤A�1.$�>ny�!��r$�x"7��K{0׊Ϗ(�x%[�i��
���nM����w^hO�M��;M�9>���c�*�ܵ���}��Z��g&������V��6�[$�L@ˆA����5��kJ��0)��)��7H��U6�v�H5�7q����L�4�K(�R���YPN��3�Uа�p���xU��r��ܓ�!R�j�Gй���J�$E*f�=:�M;3����@Ղ&:��M�XNC�:AqÿۼoњPU��9D�~m�8�l��zc׺����Ջgu0��K�H9Gx�#�4�������Wk\En��4%Fs�~�\�/�~��b�n_lU���>WC���n� ���@��9������z��ԠA�Q��d�LY������쾅�����1~��zU7p�(����Sc�7B�&��O����â�<�����ꌊ3+�?[O`�`q��Uv�ai��lw�M��M�5T�
�}i0�ڠ���U�y��hp����ə��2��E��*l�B�!omg`�� �-2�k-���J_��Fۈ�����;�#��oi��u56��,��T���R�f��/�mP�i?������8>�� H�BF�<��9�.��(ղ�A��Y���\eޠ�~?�g�+zm�<A@ڝ�Z��b�&y�&��U��G��j"撍|_-��#ge~���F"J�bW�[��/���Ķn
�f7L����y�����H�ѳﰨ?�0�.\�}9T�U0�͒�ऊ\��7y����
b�\zN$���Y��N� ��y{ ���{J�'�#�ve[]t&-ؼK��Ե�I>n�Zk:0���$t(�N���ؙ��|����'���E�E'��=n��>4ײy)�h�-#�=V.�J��zdp��֭L��AM�iJ��fH����� n�������C���VL!< 4d����{�J�Y�^�O3�s���y	㐠�d��u*�n�����~G¹��g/^�_*Nk��X6��2�@��"A_uf㪾E�F�)79�js=(�?�+����[����(3�N�YG�Gw�P��6u�*��>�ʚ�'כB�'g�M�W4~	�\䎸�_�ˎ,yEa@�|7�ْV�,p%�.�y5�,.�Q�w�OJ�6k�v�&3�� � ̓]&�oA�f>��~L,/����)s��P�����z�c�D"���Ib,K~0��jY4(f�n�K��a�(/5������?�;���Nb�o�p�o�v�X��8��t�R� �*�4h��Ҹ��l�"̳Fw�J8p�mc4`j�DC6�� ���ӫ	�q���@=�N�v�˺���9��i�=��-����w���U�m���57�0���%"���w��o�Ê=(������ �N���k�;:UϥI
ҁDCK!8�7ռ��e.�>�,���bpl�ɣ�X�`�[^r��v�/q~��8�	�0D�M�H��|�.)���V�Fwd����"
֋�B~cd?����i*I�,��n�k�5��M�
6���+����ե��v��-;���F���j�2�6Xx�U��S�S���E�dy��X��YB��&�P�rK�8N^}��{̝�b
����-&���4�K��	Q@�0 ҎO���bhJ����5kЧ� v�m=�ѷ��e�2���:X�6O�.�J�.�o*��Imt��:^���m�}.2��� �����
�iqn|����xA�5&�҈���K=P�۞/���m��,5(c�����s��lo�h���n��fw�"D����g�1�v��>+Q7`���������q��1��Ru!�Y�v��*�`�(f�I޽`��0�0�������8��OvH�pp X�T<���&ixGyj�ړq��5�Zʧy�5�U��up!�,��Z�����X\�eC'��'��")�7"JS�q���2��Q�w'&�;�{U����H���u4J�m��v��_��dO����	-gF��Q�d�8J��8!�$m�������T��g�lf_A�����0�G�	)��yDps�i���o��G����C��u��Й����0��qd��XZ-��'����vT{��jk��K�#	�
�g�NHs+A��Ԭt���֪�2 �E	�-�5���%�u�
?���K�J�߼��HEO�&��v�F2QN�F3{JdB�9��!	��{��S�1!Y��g�C۞)�8����q�Ds)���� �_���6���T�`Ӌ�����&c=#W�@j��Õ�.�F�|�"��]��8i'�l������0�,S�9R�����%�Yw�ԏa0+��Fvb��:dN@��ŋlG�䐧i�1�9�> pT-���'����g�N}�g�]�5���:���t�?7�ञF�;(;h:���$��0����tUj�Sk����-]P1DJd?�4a)Ё��'w��f�K���4/`�#�`�/���e.@�OZʗj��q�E�E�?&�qŌl�k�ľ�n:�.�C׽0���\��� ���^cw�@2A
÷�$�,��~�Z����˜@B�xo��3�6��
�����7-j�pܴb"��U�W�@���C3�$��p&���D�m%s�Z�Z˦�_(����_�Ǯ�uF�D�ݳ�rtN�!�_�e�`3�e�>�ٜn��P/��4Sg$-&�5	���q|�u�F��?g�^�ŸF�5�a�թ�?ԯWz'|������\���V�9g���c�U�B�0��"!:V�1�w����my�q�|���)ן������3�L���L�8�K�7���z*4pz��;m���V�c� ���)�9<tG���}�L���L�'�ݴ�?� ��z�����g��]IGw�T3�C�hߥ�n����C��@J��ڃ�O����#�}��ȧ�@�]�14v�k2�r'���{�T9���x�(�8ͯH�c��cm��f�m��3�P��k�>KC�W��gI�p�.F�] -��p\>R]�4O��a�s^,>�U�[��߱��R�Mm��	�p��O��!�ld�w���	�˰���q���&���;:ځNr4 �-q��R�2I�ɋ/@�}$���t`pדּ>�~?^'/���~�(��$HXZ&"��{�%��茶a�K�����t����a!��<|𯛮�`�6��?r���в�s9�1�Yi�3��&����h�(q���sh՗���kZ.�A]��z�t|L�.�5�P'�o���[���g����3��+�j�3P'9�䛱[��~��x]>�'.L�EFC�S����{8���ca�Bg��j
��B^JV�)!�zM��G��)�9��Y��>�]�~B�KE��8.m���� �eC.ۄ�Hd�-*��:FHǍ[/�_�70�gg��@�����I�gBh6[],����r}������^��F/54o�o��y([c�5�*p��5��	�>2����M�����y��e�5���
���#+F��UA�����4{����}��3A����T.��kȌD]sXU�t��2��G��H���!.M�w>����_�V=%9�I���~��
s�=?i�s&1��OA����K������K%w�ۊ�=�6zN��P��C�]��Ǵ��:~[tZ�.���9���|P�Z`�j��T%2 7��~�?���^��뵬�hޔ*��_���y��0�2�,`,$�TS�x�:D������U�&n�x9½�	�sԾJ���]R��C�������A���_�_a<�5�U�����{�������bI�U�WI��G�$��#N�Y��oX.b2Z������,�X�l��0}0:�ߺd��.SH�Z^D��������LY�s1F���[b�bѹb>O����o����l4��wn��{������\wl�UJK3up��7��M�m��az��OZ�qAl�+�/��7��S��XU�o�B8����~2�F�2@/zIAN��@����d�hF����d��\ɮ��#e1R���7L�xYh1"hevVu~��M��rm���|)�����	�{�X{��O���`�g��u�גhx�ST��D+Q��{y�I��qd�r�Q/� F��|Z���<@��f�S�Ɓ�:[�w0�U�:��s{�rle����\�r�Ҏ�Ae";���˷�Z���pݫ�U�Z�@�$�X+nU����B��T�Y'��̉^O�\Hǰ�\�P ��ƕ|ф�U�2yTI��9&X����O�_�0�!�ձ�y��-c�9~S�qT�1G����5��`7�?��R��}���?���w�%�'&[���ϫ
s��
f�:�k�u�'�EA������s�D�Xi?7SF>@sa����cK0nCF���:��t�$f.hI��^����b���ھl�ːA��Y��x"�,���(��՘�E�>Q�PW+v`�
��G
pB�e�#����3�<����d�n]���x��BɃ%R��kl��8�a�DQ�]���rE�u���QQ-q�ֆ��2F�m�$��en�̓5�a�x�p��6q;c��5�Uk�9���ln��6�΄���/�>^b�Á�>���h��1?nV���[`#
^U^X�4���B��>l3�0e�Q��Yl�s��~{�`�_��R"�3B�F��ɽ�
�Uh�O�D���Y���(�`�ݡ y�~���fKW�hts�z,�c+l�̥y��<��bHD�~;���W�euą�}&X�DmE�~�;�Z3'þ����KikcV]�_��{���k�������6B���1�!��a�4��e1�ʐ�.ב�Ň{����^��$��
��q)B������$q��%.��5\���޷*�Zyg�
�|p`q�DC����F�/o`~��U3����78�قQ��^���iL�kr덞����k�H3{�=v��k�w ��b�N��J�Ic=��U�Zl҂��A�a��ĆkW����`���33�j�V7Be-��(U�`Q�\#�����{�fJ"u
���H��]��V��_�A.�&��=�J9���~M>�e�P%�#�_8�%p�iCp�o[
���r��M95�^�`�E���:��Sô��x��@7>7��C�-!�T�����to5��
���@��0�ƍ�FZ?��]Y�J|�#�X���́���/���~���2X���0���uVz����(���ܶ�0|�E������ԳRdK(*�,Dߜ{萧]͢(v4s�y�:X���X�!���5���������5� )�q\��2�˻[t1K�
D1n��|��ST���e����Ĝ3q?,��(&9����|s��S�{v^�j�V6rZ ���:�����-��立���s�@MUY"���<�����&&�<�B ��&��0v��AJq�J�fcVrZycJϮQ�����=��H>��>D�~"Fz��Q� �t��Г���D��/&�Թe���[�%e�|�³�	䭴v˵A�A+��_����j�\����k�b�D�63l��4��O���ت�Z�^�u��Rױ~~8w�a�����,��a����$p�6 �|y�?B���1Y��y����0�Gݹh�;[ ����.��-:m��Eè��-g�>�g�jO����W��;��u��͒���m�?BP5�i����e.:JL�Ě�Y��)rk�6:Q�?���sS��,G�=�x��&�{�3�eԟN)��.��4��K�驵A�N.���(F�A"T����ZE"�"���b���o/_�J��. 1S��U����@����#�͕��Ud^N؆�Ze�P:�TQ�Qn�y#�b�-��������9��$Cu#y�c��+e.>���rb�������)Õ���j)�H��5��ź�^������GQ�rڙ��\8ِ�� n�W��d�ܜ���%�*F��̊&��T۸B
<V��Y���;�E	Q�+��W�^s�4_�teC(N%�l��� �B 0հ��-�l�Tc=��r
M#��B��dXL!���ۏt��!'�_:��x
�dT��5�O�]l���
��f�� D�<���c�
/p޺ׅR�Օv�2��6�!&�i�ȶ���#�A�w놾^��;�V�sj��o��8]nvL�쪑�b��˜���)��\�N�� ��c� y�܃���FJ��ڪ�΅��N�� �r�� ��vd��1��Z����s5RZ�?{�����4�s��c2�ϫ;�o�߬3x������^����)_@�ɽm]z���}�T����	�+���u�m���ӿ	�Đ5�#��&�)���5�8W;����v8�RI W�"[·p}�kD���������A<��l�� )����TEԩ�ś_/����沀3+o1#.Ö�YD$RV�'�d�&�[�u���)^���I�¬!wav���4S��	WD����s�<f��6�g�@��ٻ��f�N9�K7��9 ��XZ��R�K�N�.�l��eÁ{)������ly��wFWa�ވ�N����t�֑�:�CC�H�G,ߛp+�bn�sY3��TAq*2��;|a2�w�ш ɬYs꫅@�����I��T�8�5�1_J��l���$��J�g\{1o�p�IgΈ����#YԞ��T��j� %O+�vc��_%&�����a�8�*2'��%�����O��GߛYg}�U���Z�_� �G���9"#iV���B���Uࡆ$j��^`���>9�<g����Bd��I��7�ףl�M�h�9&?����� 
�#���5��d�y�'�}\X'�$��M�Nş��;e�Mcb��$*�\��Ӧa9�K�#�L ;KR�"��������+���樍�nm�_,�����(3e���]+>�,����pϒ�{('W��Ź?��R�NE�J9K�s :�m�c��V���Q�r����wHoF�?�_:�0~��|�m�P�h�� � ��C�Ʀ����aZ�Z�u��P��;�a_��ʈw�����<��omS��ݢ�N�K�������>[�$'�ɜ���mQd����v�>]
�X-�p+��d�:������S�^�K�§6�����DV�I��C�����6 �����n���*\��C��Ҳ��k{.GүR~�����B,����fҡ$���=�c��F��o�%�s5���Q1į���CVL�M�Y58��e�#�ԝ���1��W A-�u�.�`���]�i;������w��
��.���/��i� 	��vM�S�:l*K���c���*�-5s��9��/��r���'WIwR���X~aB�7��^�AA��H�*��:�~}����2b˄�T՚ր��ﱮn�B�e��U�ώ���m�$��#��X�L��w4�6Ø�'Ж�A��A}��w=�-� ̔[�pt�$��`٭t��M^����06A��i�ઇw��>��i�K/�J����N;�(��G��NF�7)�u��փ�qh�*��q�	J��A��o�Yy ��~�|��u�x߭d���#w���j�����|	��څ3�1�6���xЕ1=�d�&^��Ύ�<�}Q'a�"�a��2s6e���n�޸ѿ\���ŽpR�-�u�R�9����������ƀf�K�,l�<_��R�;h�z.U�C����n\����?�Li��D��� �k	���<L�@-U�~5�����F�7���ug�Qi�t��S�t�Ӟ9Iv�=Ό-Y���{$��!%-� ̺�|%�3�aU�N M�j,Hg�B*~���
p1$i 7�?B�!���g�OZeK�Z-t�����^ٴ��jh�>[(�:� �®*�f%�E"J�ğ���?�\cI��Έ��],�G%V?h�S�V(���)�����x�#HNW�'��9s�����0��R�_a�p��w�E��W�{k[���԰�j�n���z��Ck(P���Z�l����*E��UH�
�c	�k�G�02?���Z��T롣��Y�z��x�a��D?��*�w��m�#����T�S��o�b�8�MV�?t���V���lf�H��� G�{C�hm�� ��m@hď��e'�q������*L���-=mQ�e,}<�s����1�-^����a���)��P��*���[_�Y3������xg�0����mm�k�zG��}q	�f��C14LB���bS|G�M����׌#��@��=fV!Ԋ��i�Z�KT�3_m�y7ٺ��ه]��|�Dk���,�n2�Ș �Q9�^�D^��Z�m�D(e�M����dd��H��jl�y��`W��Pk)�cq�c!ӈ/����k�a>w��	M"��s
싉�k��z�;}��:+�Zm��~�Q���]���42��i�E��w�`�؉%*^��ZP��#��}�IpwQ_� c\k݀$ֺ���)�3|k��sX��]���p�ќ	�k0<�����h��<�x9����������\�O
�[W��Y��,�����X�r��-�O�<�e9L<��!���p&��3�	�Y������ˏ�i��?��(�]���{z4�Փا�7/�<.�3��B�wԨ��*0=V�Z�W��7�zZh��E����!��&$,�Lc1N �)�����8b�`����7v��\�����?1��bA9�۷f��&�b��6�l��ɖ9 ?��Y�俻q5�0�`ea�k�Mq]���hc�ߋ���|��X�`�z*Z����;`0#T��{'T�-�Ip��ǫ��tO�)fV�ڝ���0
�:��Ȱs�;3z���И/誚=D�H�1��} �1HʱP����&��-�Xx�3�P���Q���ޢ%[^ A6ݾ���(�R�.)nɨ�c�c
�3�(u{~�8�,GE�EN-p�#{�q������,A(���5�� ��Y�ru!!��.-$̪�����a;li!ճv�QZ�{���!�ݨ�_���KЪ2w쪔�R�h��䣠c&�\\!N���>^���Tu�)�	��2����XB�&��3//H*ݟ�J�?��wo_���I*+��\%Ѥ���ɛs��>A�+�gn��4~��
&�f���`n:��<"���7,a�7�x�zVE���I�
���ZIf:%u��t�L�����p����Fw����~P�B�;"-,@��U1�eTY��{'?��H,#��T���M~ʷ'�Ќ��K��3G=��)�s�q,�=��Yw�����b ��g���ӋߧŌ0^��!��	�cS"��|P�ǂ�k���z�S[���E�״���c��Gl����3����$ ��k�M��pWT")H��5�2�(|�^���vО�������lv"{����xJ�Ӗq�V����%�uni@��)g(Ĥ+�?|.QnbXşl=�u�<���[�~���W�r�Ƭ�l�mtz)w��~ЅT��o`�Y]�hα����Z���!������w"Nt	6�H(i��Zf��|>�S`�>8����>������Q�V&!Ce3�������X�Ɯ	��)5��^���	0!�D�����)hc�T�9蝰~"�f��d�X�h�a:��Z���2jQ`�s'p6�}�	��K�޵�º�ap6�L"��j3uZ���f����yqe���[�N������ƚ	��)�d524Z�ԷeTҒ��G^��߶K��P�<4�	6�K�~��	[:�i{��gG��U��+�<d�Ya�W��s"��^ün|���+K��}e߻��"Q#n�s�s�%�p��c0�ل�a�7!(Sl�쾩�j:/m�� �~��)bF�L4���R}1�}p���F��1ؓ~jj�z��q��/�]����Ƣ�O�u�B��&�=(dgA�*���BLT:&O�:�I��5���K�����D�xw���nJ�7J��,ӿ�I�o�(9��[�ʌ|%�����9�?��iQ$�d��S"�i���a$#VPc3�l�ے��$��X��i	��K8G�)B�Wm�;O�^��Q�H��|��hH&���Ca��|_�J��(��ə*��*��m�zjcy�,G5h��a���	��N8s�VS����D�xb_D�}<�ZπE�TXaj!j�nYŔ��y�%�3x2Q�t��j-
hʕ�u2M�mkZ�q��;��h�؋� ��?y5��S��n'��D� �PhIO�AG�3G�L�z�\rSt-Uo��%�k�XS�y�&x�W�͓�d��{&b��O;��G$�e�[�'C�i�͆��Ԑ��3�3॑ sɖ��1q�����%nqݧ'��¢-O�_͟ �ynn ��.���
)'�l�|B�:��X[�xu�=W9aX�}�&�X���k��ۏ��KT���{
{r�\�����1C�Y��n9����=�#�؉aJ�e�׋�304�T�Β�i4V!�Y�ؒNE�kA�<;�����9y�3��̀��v��S9��/��l�צ��gq����~��<7ҍ���esy������34`H���橹�{��8��J���P5�2?��Jm�}/�lc}5Eo���8ne\[+b8�I�E�O�6x)_��Zp��'@�f?	(�))=�`��������P��g�X�zF}3�<�2T6�.���p�?�ef��\�L����΀����#.�ɪ��B�S�	7��]�qG��������	�)i�\��)|�.��6�Ŗ3Gx�/[,�ցS�>�M�Fja;v�ø���{|A4�/e'�L�6&�N���I���Ia�YB��c�/ˋB�|Y��x�klT���	}hJ�x5x�Y)����uuĔS{u�ͽ�M�H��3�m�]s�r�;Yd�����)��*c��Ts�Ձ5�8!�܏ϾJ<Ҧ��6ic�լU�6���s��:+�뇜g��Y�k�*�l���u_�J���j�`��Y�/�ᚺC��f(���5����
*U����;O����g|(��X��U��]޳d5�#�][��ڷ݌#=�M��#� ���`r��n��c��v�}�^rD;���@�{��=v�|MK������X�ō�@g.F�\%a>�U���.����� `�94q�b^`ᐥ����}4̜��(Ѡ�2�03��}V%0G�K��M/���)�0��> '�~>m�6t� �ˌn�K��',�cn?95Uk�B�H6X�����!$C�Ѓ�7��db<`U�=h>�Z��p�@84�IAG�ֱW�/�F>�h�a�[�|�ҝw@	�'I�ο]���� ���N�x'�W����tp�'�n�ق�	G�'1@i��/&�C��+�;�3P��]P�u5��}�*]r�W ���L��]��R"�S�q�Rp�@���.b5�,�������6�IlW�����Lvu��/d!����J#B|6�W*mq(d�����$��s3��A������d�/�w{�\8��: �����ƜkJi�q�I�~}D���GF����h[����1��j��`�u�`l���{�8^��+@��^T����<tw`�?������<��G`HdO�Jn.�|g�_$2��)����٠x��pr����.�|���c��ߥ��<|m�U�+kCv^�X�E�e����
����	��GUh�L��R��ҏ�c��N���ܽHuE	FH�i�q��!���
�- �|�A�M�rnw��a���-��3Ċ2JWef }��CK��� >��D��,GH�I���g��W�F��ȉM$=[aM�Ǚ��{���~7�����Hq�+`������f���	�
>�HB�a�@�<�ˬ��ȡve�6i�
`e���<u7��^�v ��F=!�J���0d�Qp�C�ٿ��֬~9�3��s|(��k=�X�ڡ�+#^y�B�pQ�L���$òuO�lC��Lx5�_�0bT�"�B��َ`V�<�4CXG�v7w���Y�m�$J|�V����yY�V��j�׸o�Ȃ��F�ZD��3D�f�ƚy��}`~���S��A��ȇjDi�Y'!��k�vtۮ2�S� ���P��n���g.���S����l�,j:;c�q1m��7�i�.12�~h���;��y/gE�/��IBmG��Y��T-�^\�T����n械lFo�g�-��t�!�B�=ą����`�ݍ�MS�A��ДY���y #6���G�(�ϭ^vI�d샺g\�2jk?6�b=�^
�m�����^1��3gOK���=�-S3s"�����6H��byz:�3Ȁ�-�N�g��p}�l�K��̍�B>�g��d ��	��v���y�2t�|�n�§I��V��0��A'��w�q�Gk���$dp��7h¼eT��"�ʯ�������4�D	S7��	�~�s<�䰮�br-�@6��}J$��<�}�g�"rR��{tlo������C��-Q�K[$%����6Krlu[)/[� ��h�N''ŗ�*�o(k���������b2����0�r�f8�û�7#�*��4)���ӄ���4@�3��%�9P��ɜ~�P��E�(EAu�(�y�^��/��[}ϫ������ �X3�b��X	��J�Q�Sή��V{ǉ绖0굮槾�h�ݕ��6�/�_����&J�*�`�ĎwK��,Y,��f��j�������q�y�wi���+����
�u���4>
���:M�� |�"�*���v�h	Z>F��T���epS�&��Ϳ�'
^�q}*Q��G�6O��)��xc�b�
w'Q1�(���Shӆ토�,�_���P�k��n�j�xTR['B=3��Ky��D<��[hG�(Ō%��jO�
�t��%e�-�?MN�e��j�0'_���͌�������J�u(	W0Du�XMm�j,���:�*������ZN�;�$\��v��3����R��<=.K������L�rn��?®�v�vt�YS���r���Q3;J��5��3�ol����t� �^��D�����K��	�/}��<Ƒ{Q��&���0� v��������Q3k`�b�A��҃�T{�����rX��ᥱGj��n�9�*.?8��[��6��]ʮ.n��
o��I*�niL�bi�~`��s2�([U�Qb_`�Θ��Uκ����q�Np�?�yJ����6��$�̒T:A<Ts"?Np�`d3*� w����� WB�d78�Ib\�׳���S�d����Z#у�,�p)��j<��*?_����i1��y���b�9��O��[ t#.��JT�޿�(�����d\և^\�~���yu�*O��Bm&hl�$�r���(tsj`�u�����]�x�&��(���}�1ڳ�p�"Vr��|0]�:���s(��H
"4Rc�9tB�Tog~F:˧��i*��B��b���Y������QJ�"�L��t��`]��U����!'�R���cc1�K���)���[��L�M}|�=�54�~T�,ɕ������D��E#�����#|���rTp��7�m��'x��(cp,���x�\�6��Q�-�R�p��22�u�����&Νs�|���07���\N}}�������,=���a�g�u�&��V}'w	�/�� U:�t5�/�lԢ��"��o'6���P��%�ݔ����aO�h��\w@��@�Y��ֆ���P�W~���%7��N��0���=>&��|?J��N��ѭ0UՓ����y���4����T�)!e�w Q,�8�z_kG��gyg��_$�i֓Dѝ!o-��H�z���R����ar� )]+AI��b=�Ж�ЇT�yۦa!��ndu��L�m��
�9$�Æ�im�1���b5{�%��T��WwRk@U��V�l۳]q�rϞA���'�\�Y+#b �v;+7SzS��D���'n�\_��Q�����4D^��J���T?b�f����1�� $۔]g���x?�h�'��ь}]��?v���wV�dژ��rےֲ��IĜ{��  Q�~|Kzc���;��l�0���� <[�dC'v�Nq0�Q�KB-�/f&��iմ��ީ;g%XQo���&�	z�he�V��F��M[j�� ͨJ(<�3�T��VLKX`"�� �Ι�N7''���xA���3����@�@$�����|ZW�GPO�b��*�֗��됗�QW���.yl�k�1�)�c��Je�7&�%�c�I�����<�裟��`�����F��MP��C�lJŴ����xς�I�l�f�>m���Ɂvb�D���;GaU�{՗lI/7}��¿�� ����`��ħze�hv���<q���*4���A����HwU�H��
��*�%��r/�����@l� U񙷏����ri�a�W�~�=MR���st����8��I���\�U)���8F�X�W�n~ �Y^� KCP����a�F[�b�ͽy�Qٵ_jH�g3.��$>���:���͂cl�����b\�"��I�b �Vz�Q��s
v��0ݗ��i�ʦA�[���̗�[�eM �k��	��TεA����_���r�}C��Zc��Z���1Kе6�[��3+���;��;- İ�~7L}P�ҡv;�8�(JP�O������쬲����Uea��K�<Ql!��2
x �̺����h�@�p�Y����Kz�:!~���+��GcV5o܋ R�ax�CA���+�x���WU���o
�=��mhx\�j���t�("%��\��9�PN�Q��'��61�-ŀ�qW
�K��8t�˿e�{Eӎ�r��'��&�K�6�E��raw�I���3J,ć ��z�����,i�4YT��M̫qbU���)��`�:N���}Ӝ?n͢.`#���i2���<J����J�ZÄt�_��i������N�l\_�s��&�Y��z�=����+^d"��R�K����<u�XU�;j7���5v�e�A��Gݟ�}:���B���c�Fo�Hxl�wny���/�'5��Q��ԑk<k�{X5T�P��-�c'(u�Q�#�z-�ħ�%6�=����?i>�FaBW�Sj�tt����f��l"���Y�j�ǮeI^+�+���a�zP^�~�NƖ��Fq��|�:<]�תp�T�b_�f4�W�n"`��1(,L�x�U�v����,���i�O�{�$���i��	ou��x��]s��!c��K���8����_$���S0M�: ��pgm庼!�f��`$��m]i�=�
�|�F���Z�Nz��K)�F3��m@�H�����>��x�z���8�a���H;��/�2�ݸ����h`~��;|�ƽT�/y�,xK �_x%��삧0^��8�&hC�ګ�4ҝ}L�'�bcy�:!�H���j�0�Qd��7z�;�^�Ԋ��W����xj��JD�":{JމË(�2�=._�u�&�L�,ӽT�5s��SB��v�(m�,���Ȯ;">��CoŠ9� Jf�o����|I_�y^�5���i-�Sy'�Z�
��ѾǑ�~�O��A哬�7��@��!U���e&w�9&8	'%�V�ޏi�֠��c�',(5)h�X	�T	���DH��pJ��Z��*r�2��� �����_>���<���()<[YI�Gt�l�X��9F�eurv��}>O��uQ���ysO^'/��aW�G��+c
�I�:~����?Z֦�N��xJQ��|������]���)]���[�>�0x�&,7߱�8�=ǝ�Jʓ�~y�wKC|B���Ohj��D��e�s`Aw���v~�yqJ1�2�&zp��^�c�o��GJ��ud�Kf��SD�q3R��{���D�?*�ɇ�g)����(T��;<%�忢�P~��~j�U�L��zK��z�81z��!�6�����ґ	�(�S�y=}�҄h;w����V,[�dR�V���7/C���^핵w[��	4����4���u@Ӵ��T���!	^��X\�
6Ha�gP�lit l?�n��T��|��2�=�OHO��T�Rcr���!Z�������s�X-�z��9$7	��<*����1Sysã��#����.K����ؓ�����$�oG.f$u�^��M�5����_D���IQ�	�#���9�M��u9ا��)�!E�K���)³2�[-'� Qufl"P�u#��ʌ�T�1��	+�ED]tc�vm� X��.���r��E�����)�\�i���1�2R	��&6,n;@I�U��Q��R)N/j�ī�,�fXFV��>�(xU��K�*���M�အ����Z�������OU�Tl�N�V��X�j�q����Bt�c�#�p�!,�$�I.gE����gD�9Z�0���@�:,�i���uZy��W7.T�S`^��Jj�ԧ�s��4��NN��SӍ>�� �	;�$�V@:�h]N�`IHG�D��5�虚���'9M�n�ZldO�O��>���H0;YZ�*ӱ_l4A�8~F�,�Dp)�w�!�_�|��m�c��M?�n��������b�e�:B80��L�xg�dx~Ԝ�w7��'1��^�a:��y'��&q2�G��!΀�����؃gꊧ�8�Ϩ�]���Ho�f���h�9�Sʠ:5a�廉n.�п�_5n��~�?z���6ѷ-�c<��Ԣ2��j싪��5�BAP�G�GkʜD.��/^�>,�Y:�2He;�R����]���z'#O��(����hv�'�r*y�6� w��&Z�� �w�^*��c�py���}��I]��N�÷����]f��?窂�8Xv��vy����,R���R�}�U��;aBPazp[�� �pl̞�~�i��<�i��f��uN���q����H�~Żۡ�	ؕڪ
�'U�P*��o%�@)ۀ��[�⢆���<J�"���=̬��qc��T�vv���B��}�0�7������\RBG�'�[X�a��b�@5�s�!>#��B��ԏX=YB������iE֚�u��+�Y�rI�����;�`�iZ>Ͳ��Y�`d� �5�Ҩ���U�{-��/~�.��<~'�r{i��`D`���{h�h�E`�e��t�|n�.9�M@h�~#f���)�
�̣���$�t^@?�T�Z��7�:ܖ��v^ų���l�e�NMo~�2�=�偩����Ƒ���^�툃xA��6�=�	[�����Q��M�0������$��n�Ux��ěo �^І�>Cv�3�
���Δ��]ݷу�rkM)R�kF����t�肻,4�p�ay	� ��Y'|E�ɇ _sl���S;�|qg���מr+n����?��Ї �
�SXu���
�$"� K��6P����'�_Ŭ~�j�H�_�vs~��36\�柲دZ��@{վ,�$>@*l�c�:Qrl���@�u��T\�3��*����0�ci�{Mqt�zL���l�����T`��w�VȢ�G�>��܄¶;>����BB�r݅�c{�]��^hhT��d�3S{-\�!�IU$0���)��M�0܂c.�B�)���+�/o��^_x���&��3�Mg�"��4��k^�X���o�h7O�Y.��m�og�j�F�X���a�-,-]�ZE&[���zORu�5��|��$gީ�t�5�V����Q�����)��PC���"F��Su��T9��n]�57U�hy��8GZ�����<��_�'�b�39rb	�Η���r���ܟ��t֮�Vw�k���U`ׅ��y���a�K�!���Y�,o?�\� 8�i�����
�Ģ�����Ň'�"99Q�V��)�4H�f %@w���2ə�qq[�(�Ld>m� O��)�q���$�z�$^Ƒ���Z�V�~&���>��x��?��fCQAKY�R]"E���'Rg���6U��Y{.f"��A��#�}�,RWgc����ZW�y��NVP���,�����Ƌ��u��{��^���,|j���`�^dm$ ��$��|���QQȣ~���{'_C��D�U����e�B��#�̔�b'G�k���=I��(��IJ"O�[��OF���KB����-W��@�[ON��\-l�����R��ָ��Z�b���a�T���-��sE���p��~�@�SYD0s��s���ǡ8��\q�lA�*�����,���n�k�ikC_m���<���~�"ձ�[�&���1 @DK�kcGBsmet�ܶv�Ӧ@��X�)��k:;8ȕ�^U���;�ӧ�!��T�	��{h�H�@0CX�Ad�w�F��|�-�B��mA6�߰�1�"{�$�z��[q�d%/<�	�\�N�ǸE;�5ћ�������l�AI��%�V�U�;�~I|����?a�|�2��+4�x�����}tʱb:ITd2�;$�g��9X���x�@���|�~�`
���}��'x�T����j��#��ˀ?F����5��+�#^[#����k�mĺ�7̡b��^.����ь���so=�d��r�]?CwB��-����e."�*�lF[ߊ��h��(_tz)�uE�?"�{m!2�|%�s��X#�S�ҹ�?b�\��)�$"�O���O���0,�4�9{�*Vg�Ց�ڎMp�� mظ���$v���Q�״
?��Ӽ�}�Go�(��N��̀߂K������H��~\�Y[��k88�7��G��"���b{�rK3���$���#Y�i!������LK'��
q��n�[��Bz��@=�Χ�f���9�FP����Ky��`��ܶ����e9��]Ut߬��:�{� ����/��lb��7�� ^d�%hHҤ硜��ZAHK�_-EXs]����
`U��Gq|X/�^b̳�s윒��4�ˮaK�U�aR	Ȳ�
<�uv�����!�-���S���/��|CS�l �ڬx�3��N-0���lg���e6_�ftօ3!d;�b����	�l���[r_*QfH~nX�3��Y��da���kk���ǜscO��_W�fx���/$ ��!^�|����:�	;�=Uj�R�|�؋*/�I�D�-Q�"�=R3v�%s�c�R�����Ƽ�-�����߂_ii�s�6~wg�g�)��.��A�� �Z�7�Q�Q�|�������룳��(��7�.�a�~{�.�Ǆ.�����;ɊV9����=(\�j�<p#:	����>���ge[;�_y��R�E�����Į�}g��c�3�u?O&���e�H�$v?�[��E�o�<<�o�G����d:�Q�%����^n�\n��T��-/,#�m+�:3^�/S�^)'��>�����ۉ(t_֩Dr��$웻�5�ug�;����X�o�.�C	��H����h� � ���W�Ȉg9~�
*�U%�T�v����})���6~>_Q�S>K �&�Q�Q0�� Y�6��E(����ǎ��eq�9���@�ԁ9��-I�$eo����Uq�HܡP�'���&���$^5$���e��3T�c�8J���,�%ű�Q������%�x'fj㽘Q������V3%��/3���,�\������{P�gze����m�����9������W�I��u͘S�)i��;�w ����#*+����N"/(3N��C-��C��|��cZ���4��Aa�-�[_]�GH����%ד����<���������?��왖*�ϝ���4f`�k���0rt�	�H
�j��@oI�{�O��{���av7�TPe�؅���Ʀc��^e]�V�B
�H$������.�f��yc��U�|��c.�	��6�U�(��|[�`����G�������h�va�d�&4k_b���j�ҷ�b��T�Q����M�D�W)��BI�%�9��g�̭9G���hRD%4��-)	Q������� �%��$�3ޯl~J�H`���B�d@���_&L�f�l��Cx,
dvvb�����c��e,(:��_�����BE�=K������9�#�;�eF����=��ɨ��׻��4�.�l����q�1Q�8%#jQ��b�}���IAJ��ϲ|)V���}����Z`�;� ��W�/]a�*��~sF	�Ľ@EԲe�C��j�ڷ��v�H<�;�Ο�3,3�qn�z+�^N?���ˠ��no`�7�޻0�koťD�2.�=�\d�qW�x��Ԡ�C�w����+Q�*��ߙkG�a��Wk����N^��3�Wnc<���l+���᫐�M�q��4�����:U�?�C�J�kA"��Ī�^���<g���
#�ox��xx$Ckw�!�L}�w�ɕ�8�=��S_�{�f�k0���H���q*����v�%1�	���)�z��Fz�9����s�4K��U(�.vt���	/q����LCP�E
}WG�2�N�Y `u�|5?�����;7kDY�C��dj��A��d).B��u,��^4R�hLs[8y+2�/��6��-J�-.��΍��v���]g(�Xå��DXi@��$5��*E2_���|����W�ZQ�JD��u��GW�
5 ē�7E�B�s2_g�����3Mz�?�˦�\��*gY2 ��c�O9�a��i�GL��:ȇ3���i���Â���� ��g���<l�폤όC4��_����W�z+��������9{�ndwb4�ov�Ib3�3�q53�O�lK�*J�4��%�s��Xiw�^���`���O���|�ڋR��!�
��o�ޠ~b��XU��`��Oֹ��9�'@�:��'�Y�œY��J?��B�TQ�i��J�����"�< A����X��	F��"u��~4x�/��Ɛ�g�@|���w��.N������۵
M2u[�#@�/Ц����K��iIg2^cNO��
��޼�{�|�	�4c:�H��x�3pv��qOK�lr��U��D_{'iO�Ѳg�ף�ZBMW�cڀm��3n�Ѝ회��#T�0��U�����iD��2Zۅ�y�K�c�.wr�4���b���,��`���B��I̐Di�'x!�J"e=h�X�ƊK1Ξ����8�0'u����+�*)(Q)�����^z�Q1����b��M�Woѵ�-3��ԔPw[��D-�ڨkn3��'B��:��_5��7��9��P���� p� ���YA�4�&k+��P��$]�K�L�}ZuHx+%�����{����Ǫ����,>}�Î������U	�p���~>��`T��U�v��Hm�`�2�Xyo��k�s&��Zc�tΜ����z>l��v˥�s������؃��8wJ����4��i���yA�^Ld���-�T������1�>�w�0�X�n�xH�m�������{nXg)&���X0�?�t�"��1�k�x��#�� �l+��7�3�7qHg
ע�
~21�t�d��J�:���Vy�APԔ��"Q��ZS�@�Q���K-�ʷ�����t���*q�!617�Z?D9UF��L�|`��ʒkd����9��u�X��5��3���	w�4���sv�$̇�B��F)�O°z�0d�J$�	���u=�׍:D��t����������;���<�X$0�DM�~Q Z�W��񯀚�6�]t��
�͓[����8�pQ[-���TWL,�A~^��:
�Ǹ�E�֭fA9W
����F�K뇵`[BWl(�才;f�=�Bt�rЋ�~���i�9��y|N��b���<!��b>�{�"�/�z'�(�u�X���/bq��5g)���*��NFx�.�Y�+_B=�J|���M���4���}�:�5+��P}/�M����sv�̸<�!]�N��Q��f��	�*l_1�#�8U�B��R���Jw�J�Ċ���.Z�nX�G}E;��J�=M�~�;�5�&�h���;���.vv�?�8N��ɚ��(g�q�%	���7�\H�`�����l X�a�"�3��X�q��QeFv�9�,�儍�����}�\�]�D�,1�ѭ�_Ru����T��T�����?��(h�n���{@(vF.���o�d���%*eB@[r\�M��� ;ʌ�w�s�%��ě|
�G
3�m,�k����?D � �2:�HB����ݺYB��� U9��[�C߾
3�&r#7v,G8U!?ر[1`ewL��
��-h��<�7�y��Z�G�'��I4ɖ>7��E��)_��c5l�X^��8��N�~oڔ��{�f.�a�n8ݒ��E�\¶��å/iOܳjzg�y�\����阐8^	�����ڡ���A�i�f��!tkO���a�&�专�t�����M��1l:uLdx:i�����3�(P"�kC���YP���D���Ix��w�D-�@-�6=�6o$	��%�W�����£��� R[�GT�?D��r5o�A_�k��,476�N�D��j�W��օ����/W�������@��Ka�z�{�#j��_��F-�`���V^�.�B+ms����GsHSY��8��i���m��5���1\���܌��T��N=��BZ�D�Ϥn���j��.}��EM�\���s�R�nN�`W4U���G��.��u�?�e�P.,�)��+#���:ZG�O�Ol,��<Ns圆i8J~�!k�yႩ��a��$i��� ��z��vw�c���oK����}�l�ھkY,�'�rk�n��] �L'�s�,�#b�'m�)Ѹ�sL�-R"�����z��ᓣA��I!sz�A�����\���$�V0L��W��ka^j~\E��f���cq0IG�*��9r���Fu>�P�f��� ���z���\��6jd!}^�a~yu*�̐���Xf7d�쎍_s�v����2 FGG�w�;�w����݃��@C�0�pPy��	��M�qd7Cs�T4P�6��W��d|A!$��LW�{�k6�D-$'ri��;�K���G��`0�jw�.��9K��[�a���Nkk�y�'�:ɌV~�����I=&?_4�09J�~/�G����H۠;2��l�n@�w�ğ �]��L�#Y��]���7^�`����w�q���*1�M�0[�p�Ӕ��^݄ir<���Bz�cm�A��U'��$E�J�\:�^!�C��)��ã/�,W��X��`�]}��/{ܣ�����y��+EԜ!_�H�`F���Q���j��)��<�k��'"��p9�����<����7��.r\W��A��v���`���L���2�>����'Ή�~07�o���r��Ԟ؃Ӌ��c�)�J���}�T�.��%�)�6#T�K�CNX�S+arQ]��w�EPԷ�uH��k��	^�*[�YǕӟKl ��9�y��g�7�Lk�fW��<�t���.Z��ѧh�3�v�Vgȿ����!ʄ3�_��؍n?�z��s��ӭWE8�}:�gJ��z>�;�c�Wh��x��jj�J�TU!}���d㾤-�c܉6X�z@�ykI v���I��'~�z阆� \�նqUb�r�y��n�Hr�(��Z�7W���K��S�[;6�;^?:��7,�ӫ��hχ�U�گ,��M�9�ߓ�V@K0���Z�p���h��#�z�27��٦�:�+���x���|3$Y��y$3d=�q��$?���}o�����J��B�^8Z��n�%�`���U�
VҀ���H�G�Y�EO��35#!�M���j�%�?搛B`LOḐ�2������g:�ow����>A+��,ʝF9+o�֓�!ۉ�*$��%�&�)�*��1a�m F��n�`�e�`F��h5�(�$,���4�YH�[n�<�:�-�`H���۬&�#�ߖswƖ�������D(���]� RM������h�dUzBj�㴥����M���6IĨ�Z!�B�ho��0�4��AQꂫL�z�:�?6�G�҂�������&N<�qΛc�U �4�a33� 	�[c~.��H��M�b+�A\y���t���M�$�� b:;W:�[���>�LƎ`7�~�ל�}T��W�D>��4�Fn�&������4�A�R:'ꌞ�O�{�-��-ɟ�I�A�A0kLY�'����cj޹�=���~���N��!�ԝ����.��Ae���ι�'ޫ��b��T�<���Stk7� ��f��N:)�T�c��@��6DNN�s����yqk����;�m	S?idy�`����	n� �3Y����/���N�Nk��m�W���q�Df����E1��߃p���!b�0��|�_9I�=�0�i ���,Es�K������%˷��g�<� �	FҾ|;����[n�Y�������P��-���kn�����a^�ֱN�a������X�RWJ�2J�yS(�P/�Z0׽WG,�!B�~/����L�Rs�ċ
BYu<�]^p��$iED�:�C�Z�,������p��m�+wcF�QH�>j�M���#U���� ^L��&��b�KO�B`҈|-��ؾ]�¶P�f�X�^�Һ�v����d�E��
�٘�׿8����DC�=4]�j��=o|�S#�'cv<}�Χ������-Zn[$�E�����$��$֥�g �7~����	��X�p.�?�����k�?�ԕJWG�MM�7�]t����dM&������N~�V�Pћɫ���ý�i�HvU60֮�Ֆ�ۏ��d܅A�.s�K�ܧ�����Wz�.�Y��f�߄�o�a��A9�p��c������lC��'�v�maD��� (�R�+y����=	��sߥ
/K��Z����d&�YEC���uK���K)�Q���Y�@�ř��P�V	�l0��G>Y/`���˫wҘd����&�I9r��W�FT����8����ES�U`;�~v��h�39�����=ո��GQ��H_���ءL��h��3���C�o��q�a,S�C)��ך�q���M%�%ɳ���l"��G�;㴰����3�7�`���-9�hg��-�����3p�F�q�$}B��N��6�⫪BAT�_�s�eD=��Zt?a$I:J:5����O2GUv�Y.��W���?;�$�nm�N��m���l����N�
L��R�~;�E���W4Y�������5;܍��̼ `aZn�ZK
i7{�����5O��$
�1��˴f�3�ݺ�P(�i�ip&"��Ҁ�-��84�6�}�2qL�OwU!����P�I��#���8���l�(M݈���]�?ұC�sE�HH��E�fo�?��C�&�(��v��[y�wC�4��C�HaV�ı������'	@���q�Y3��'j�;�����e�r�*R:��U;Z?V.�x����y����k�U	
�hu}iQb�2ź�.hs����`��Ÿ&R��[����fh�&N�$��@R���}�E`C��� �f��H�P����|��	`��U.<�f����I���uq�#�i3��)8׫�	�Y~.*(鷛F:i|����k��	�S[_�d�?JO��au8B��Q#��n��<3�A�6}���#@I<<���VXbH�&q��*���E9�(�2�0�Y̔&e���f�n��똇�r��|�h���cr(���
+�HV��^t'�Wp�w�L=F�
�Ϊ�����X��
��<1e���F���N�hEl��@ dM�bE���fdT����%��)�� �� .ȅ��;U����G�A��C�[���ބ�SϨ�L�8��bcr�jg�'8�@� 4��B�>���)m�:G�˜h���8eC���n��L�r�@��ߠ�!p�[q�Tة�n<w�e|T2�b��|�F����OQ��G~٘q�I� �,�D|7��gy�ݜ������Ϳ͐2����g�L������&n�ሱ�f\z�8l�:� MHSΫS"gù0vu���y�O�1�Lq���� >�g�1:&���+�ǙE�<��>O]!��c�ޱ�3s����s*��+���׵�����< R`����g�_��2(�ؒ}j�f)6@�0����;h�T�JV{Z�Gc���wܨ��30,ZS�"������`I����4�d�	�jcP/���33�on���k�>͡'dSjt�D?��xB��{���kB��o�㔳�WgO�c'*��WS�� ��5~^��X�N5�g�}ى����Jvf/�Ǘ Ok�������=˽�)��M����35�,�)+�oO��*��C�Zg�l������*��<�Y%E���,�|2|�R^ү�$} S>�^!��5�D�r���g��%��g=Ō�����*�@����_�������c��G��D�K*�3�!�$�B:c[>eU����YW�W$j�g�گ���ܵ���Z���<�>����'��,Y@�����*��ԙ{�|}�R�.���m3T���h�8eƴ��Y2Ƈ�i�����f� U���D��9t��
�cI�"���h�'f��K�N̮z���ss3z��7�s�#S��ϛ����l :�u�ey3C��T`&���;'�`4ZF~NZ��2C�6  ��1�5�X������%0O�X�V���b���3Oc��_s�g3sL�I�␱��}��g�d*�U�a�,9��� x�z`L�ǐHf��|�W�N�\m��&:{���^'�t��q�;��Ow|�/O�J� ����ؓ�9�����$6U.�q�魱ӾV�b������_G�s�(��ƚ�geu�D��6S?�Q�N���9+��'t��b�Ϸ�:��l:91�����i �*��Y*jp��� !3�� ���ғ�4_ӹ���fɶ�Ig���%�N��A֮�1��R\i�;�Y�.1����p�/��`�g���]���1�x��N�t��[�ԽV�
澫'�&u]�g'fyDZq�`!v���a;�I��3�S�}��:���Lsk���{����b2�'>Q��Zt���v�6�cò �e��D����3h���E��@�:�:<��T*�.译��80�����M�z�kH�f�M=��x���J9�C�l`��`�%ZS���@���/���Kßz���-'�g6�隿egN�D�p�Fv��V�B�>��vC}WV�qX+}⑮Z�z��ʝ��.8R�;�!T�-5>��7���)FXXײ��/{(6T���Wv�r��%^���2����b@KJ�%ne�2S�����kH�9y�[�M�U@�z���8�5]��J�ͫ*�4�JhZ� 0Mb}(̓��-n�Sng�h���r��8�Z�(���ȉ/oa�-�R'P��T����1
�O8��7�!�1୲Y���1F�WS�3�{Bl���C��	Ir��0�Ȧ��$c� �؎#���;o���;�7�%LD�/�M��!���P|����<Ac!`��
*��d��n�VĬ�u�r��������J��!ˌ�-����%R���c����A������"��&,�ϝE�9�DJ�l﷔ҭP;��T�1��b�%�{�������fq[<Ȍ���
�A��g1y����6p�� i����������mQ~A�(-٧P
���BO��)�-Tr�^��I+�a��T�ɬ�)����G^�?kd��f�AT�7��[`�M��?�h����*nd�'����7+N��>�#�t`��/]�៎r*�U9aeveX@��%/��mǥG>rd!��Hn��w�l垆w��p�ċߦ8İ�H���R��)2 p��`a*�xlІ)QufW��XnL������?�C�b��^�Mkr�CP��c�jǏ���!�L�gK��ͪ��o&�x��คԥ��+�(�7�ٞj�/m7
/??�/�$�K6�l"x��w%v�m������X�}7���2�p}PnFub-� "5��i%�{�g�et��{�@UJ����Gb��ʝ%82�ڦ�O�__�[/��X�s2.��à��1�p�һM&�M�8m!�Ai���S�mZ4}�a��q�	���)���<tM�b!5h�;��f=}`5	�w6�77@*e�8����������}�uC���~��@A��:�������"�ڥ������[9s�ʎ&�,�*Yl�K�W���]�����+MƊ�:@{��:F�����ޤ
���n�v��n��=�d�sF?��T��O�ꇟ����N&��=y������,N-��Gk{�&�nQ���ǣD�?sPۿ<{�I�7� X�̼����`�}|�\���v�0#U����/�Xi���;qS�AC����z�#|���U��΍Þc�=q���|md-�I�
��ܑn&c���L��֙�����;'s�Zv�a�`���km4*һ���ej7Z�)��I�Y�y�C��?-�3v:E��JE����U���j�1����U�#�cAE���Br�7Hx9�ݹ�^��&c�)�X����]<����~�msD�v�P54
����{���vSd0��ӍW�26��@�N����n1�ٯ�з=|͸��w�5ߜ�ԕk3!"��D׾�|���� �S0EW�^oԤ3���X�E6��ö��5��s�Kd�xKwY�3�X�N�:*p*���ANt�#Ψ�1gIʨ�9#�sV�g;��ڟ��BC#H���ر����;[EFU�Pd�R[�_~uGk����]�w��Q�_ԳC.p�{���Vu[�칍��� 	����I�t�)��8������$^��K���'��^������.smX_Ef������qʹ	T��<,��K��}t[�/u���hr��%�� >yYgr:�я�@�.��u����ퟹ`�g�XU�:Y�����Պb�d�?�I��]�3nL���A�]�����d�]^�v]��n��U@����<Gr�MM��N����~"B�o��g��1G����NbmO�@��n:SMCZDZ�GXD�p�r|	����fQy�u�{3���7w2���%j�Ǚ�I�|�uXg%�����׭g�����a��� /��L�7\
��E(@1��D���lju0&��X��	�iB)��O���k�FM��Ol���]���x���\��4Ą\��
�C�k���%:\���S�<�b�{��B��~�F,�z:S(a`z��q6e[|��I�:u�!���r�RE]tA�t��K1e� !Al%�[�j&�N��#$P��}��-L��qs��t���\6�OJP��CΣ������!S���M�����iFVp�e8�e?�q�HB�#jP�@�E�zm�/�7��3B R<N%=���mW�o+�����Ǯ�~�������,�S��$|����,:��{���K���h>�c����m�n��w]����HnXE�d�Q����T9U���\!�/ <��,�;"cJ!3��s����P4�Mp,�0{_6�{�%{3-i�8�\<��d���Q�w O'���,���q��k�h���K�8W��wv
�pb]���D�3>���� ���b�z������W�<���l���t�Cǌ�2�d�)�a����^�`�b&�´�*j�d���M��k�d��d��f<��+��Vh��K��#�o'�:)��{�93`Vc��_27@n�^`{@1�(�םè����5L�e���A�
Y4Z�f��~3uJL�P-����7�	�X��ӯ�i����z�R��,�ʶ�����W"�+����0�1�f�tQ�c}�4P�9O10܀>�st���ϋ_g�3�ncL���xTH� ����]3�<��k��E>����_��M���q9O���cFC@6BM�`'�6�����K,x���r�f��:ݾzy����d����m��ը��l�ؘQC�9�X��39�m�,�i���A�3F4XZ��J��V'g��5�_�����Yq}�� ���=�F��x�!H�G��^";�Ex1��G�䄋�P>��.V6�RnD��y A\����ɗZ��ֹu_�o!��e����= q|��<��~�nJ��wl5�(��1���<?[!��Em��Q-�N:���Tj�o�(���%y[�"ҏq8�Pi�U�;��o�������������%�!��vK<�DP:�P\?�}m�Y�C2���.���H��h>��h�g��6�9#`�'_@�	���c�l��k��@F����kщ��^7����Sj8C�9����A��{.�ȸf؜��j����RR��M�J�'�9J��9ҽנK��X�y�M�/�(>��-C�j$�!/�乭UP���=�)u7 {r:TW�_t����3|aٸqı�iPqA��aT9���>=��$L­SEJ����tk�4K�r��X�h��0y���^��ovɮ������5f��N�*J�(�F���_9p�&qۉ����&�\uu��e�8�1=� Y��?H=���fs&�w5�#�?
�v��
a5�՗-�7���)01����1nX?gh��~�\�r�q�.vn�'G���>�l��/�:y�u��H�/��?�J�J��52/�쿬��$��Th|��
�%d�p��D�Ƃ�m3���4��Q(��+Qfg�st�����3K�O�I��h��1,����ּqZ'N8Q�k�	�>�c����"h=eB�:���5���U�&��oe� �ޡ�4�\�c���j�e�M�y9����E�+��1b���������vP��9���Ku,�Z�]�እ����^�&L��l�L��dȣ��U�"�]��)��*;��[�0�oxa-["��-2����$�ެ��������^�/}��w!����'�����O��v�(���9��4������b��'������<�'��n/�A�mN�c�&^a��AJw|RmS!�x�M� �
��{?L���#u$T��y.�~SÁ�G`��>��;Ѽ:���!5ozx)fY�J �T��r]��wz$�Zk!�pyXS��`�T&Va|ۍZ�>�%g�Ҿ�hYj���>�#�k]��s�AR��SCm�x����Z�q"W+e0��bl�9����jcD�j�F�ԟ>◗�f�R^��7�z,�i�Q��H!Vћ	�er�-/�H�7r ������{��S�y#$���i�R�ޣ�6Ƒ{�i�=9WCb�"�� ���l��	�����-���k:�ts�F¡:����)���,Ѣ!�����p�c|��c����� V��D��d;�2��;�ߵ�Y��U|+�_�������n�rf3%y��j�y6�P�"��U��]�i��~���H* ��<�����˼�in��-����K�G_����'�H��F��Bq�&-O�v���gv;�ѐ�gƛ*
�ʛ[7�9q�᧨J6ʒB�ag&�z?K�0��Bب����Đؠ݂�[_�4bA՟��B�>���^����.�I��-��һbC� g��f6���$�6�_^x��ܶ�6��j���	���7+�b�Qk$��/����i��_*I�	���J�8XS��.�M��j@�t�2ǐ��X}�nѱda"�i�5G�a���޹l�`O�5�<�]�H�+���]��1!N\�~��~Ʉ�D��E	1��23V1;q8F��A*����/��s�}�~�R�j�E�4AޯunQ�I�5b)�^�O^�l�b,{�8O"�* ��Bq$�c����7A�1?	�0	���!p�P��&΂�Lu5!4XF]�E�[4��T@�KY�sO�Iש0H�[>%JZ#����u���H�����������P%۪�ﷷ��a�C���&!0��87y�!I�������!&΂��7��ߪv�6����/�cl�
�kG��ݵ��^>�qU�+�ԒƩ���N�Z��de��9��P����LH\��^�}>*x�s�	�5�����ɻ�i������sa��Z�$`����)��M\|�'Ǭ�X���C_ȅF8���rԒ�j���z���F�$�@�k�l�`��� �� �ɘ���c��2��DESC�����3���Y}ˠ���(܏!�����E�\n�p�o:K,57�
DI:�Qs'<b&59���;����sXZ��Bu�1N_q$�\'4��G�����@�M&���D9��Nu���K��B�.�]�0~�J���L�CHl��&$=���h��E���H��Ԑ�s�v�fU~M�ׂ_����<� M�5ó^����E?�8��F�z�	���Tv(+��z�49�����%x������S���%���C����"e�9A�J �,kC'rB3��ed��!f3evmU�tp��@�-�`r"m������Rg�8X~׫w��X�c
���p��5�\�
=�����^�kV.�sJ����&�C�怾���׀i����cR��#>�EN�g!�wS��'�����k�)&>��n1�������78
97O�!�[z����Ǡ4w6�Ku,��
�3�{#�߼��^?��h�l_鼟Y� �L��^�@���rA���dl_0P����� �P&g��ф�a�ؤ'���lIbt=��`�d��d�!�_�N���5˾�P��F��HG�v�W���*�ȽB�s����K�F+Fw���6r�}�}�t������yq��Q6�R�YD��o�Q��\���uy��S��'eN���j�[�BNO]ک������q�+�3�]9")��BKlv�%Yp�m�ƌ\�����)�vY�;UɊ��_^9?\�zhG�̪����q{1�Υ��(�D�-^f|��' �SK
m�q�a{��\X�{�|t��
�tܗZ��C+c��.���G�	+�`�˹nv 4v���%>�o��MV"Bf���3G��u1r�LHi�.�p�U�4��>ZN�*{��GU�N��\������!��X4�ƚ�܄!/�Y�\��&n
�1�$9��s����$��v��9�ó��k�SȻRޤx���Fx.�U�p���o��;�7r��2�*���:�*�to`O�s+��,L���q�@�"l��$Ipm���3ڳ:�P�B���o]l~J �nk�o��ʗ�uF9���}���3]��x��?@7�%�$�I���2w�|�lʍ���@�N��]��<3����rVx�r�٨ա�$u�b�T�nـ�r<'V�O�f�8����,�i��u��`�����% )i
�~�)ո9s)|k�W�	�ʹ���l���j-����5Y3M�q�ߊRT0oF���m��I��sR!��S�X2�܉�䴕񸛓ǿU�s:� 5$�E(A�5Fl�w�i$�o�R��m�G�lS(���o��	C�j�l�)-O���z�Y�<A�i����#TV���x�+/Ќ� �$��0E�O\v$�޼�~�wgwMf� )V������B4�t�S.�´)c$"�����p�σ>��x�ߐ�;Y�ʻ3��o#�a��A]s�J�t��y5�HMu��P!`l���	D`f��.`H����Nҵ0a�?
����ǬXӍp�cE��,%Y�������}�^��8�/�������և)��6.��#��hG�V�`���:a�Gxٔ=S�����m��ܵ�N� 륱+n�SV� )���Z|�B7΍�n�;���Vmt�Q9
.�/�*�.by�h�e|4b+ ���f'YE���>���Nc�3e]s�ZJ3��_���s-�̵_��/�=��x�(��Y�p�]�1=�Q��)9� ")X�Rҟ_������c����6��#�>�-_�hS��^���Xc�.,r�Slٺ�
�(&�߰��8&x��r~_mp�ꧮN1�}��{;�"O���ݘ[z*6�����]4�q��H���"�];qiك���r�jj�<�X:,\����i��b};g����z5Z����v e���0R����ժ�����C�K�f�/����Ns���'#|�G�r��u��n�b�����td"��Q�pN�eڝ�~�Ʈt��po�>�'����Z����>m�\{p� ��9�[G[��_�?<7���8\"��1^Ni'�YK�q
���6`�W�qtވ��Ny6c(����]��{����l3�H��N�m}b!���T8f9�U��ʓ�گ�! �sH�B�?�/vO�@�j�O�2�R�4�K�q;=�ɂp��/�ₒ�v��P�-�@<�CMn�Ҙ�)y�	5ed4����y�~��Z����O�nB4z�I�?*����1}t�P瑇�%���Hq��_����R��n~�t�2��[�o���.�ޯ% ��M�}�`fh:$ݸGq�ҽzۛ�f[���s���.h�?�����0PA}��4�]����?�(zY���$���0G�LR�ʦ�	�p��W�O��Ɠ���)!��<H��~t�O�OO%-� :u#�Ӯ�t����z$`���{�:l�E�O�}�%�Wṡ���fi�����o~�4���>\4�y�����RKU�|��L�D!f�ߘv�'6>_�z�%x4���-���xM7���m2� y�x65��Bi����3�t v��T9Q�3�'<�.�n>wΧ򇪧m6�Aޖ��D��i��H=l��Q�
��A��n%�C@���?�+@>��G�<A�K�YtT���C�x�߮��P?�k�m���&{�t^&9�I~V�����s��q�\���1��L�g@%_��sm�nO�~X쉁H�!�>P���n�?��$cI;H���h�+� '���!e���y�+�jl���$C�c��&�O�c醘D&7���:r�}��K�y�-��^��Tܦ�4"���R~;;㼣���P�H-t�Q_�~&d'=JL�Ff<z�|x�)�g5�\4J��V Z^K\�V�� _�F��Ķ#9vx}�7��?h�~�ƕA>8t
�h{H�{�_�!G �H���.�����\�8o���,n�:/X��,�k�]�1q����G��q��z�Ҝ��Z\�p��f�\c�M����	���W��Y��?�=�����d z���1����LC|����7E�d{/��6�È��v�mA�e���	j��|�q��rX}�9sESs:�%�+b�y2+6&�jmd��? �;��~��kb�s�`��r� ����~(����Ȼ�f{ͣ����gR��M��Ĭͼ]<3�!cJ�S!(���ݑ�����_amm.�#���-9��(�Eߜ��ޫ��L�$�/^�%�S�P�D�����$vu�Q�H����m���ܾ+CϢ����:�G��J�t�lk� f��*�~u����)�,?�e0+M��8o+S��ߕA$](�dv���L��t�7���@Xk����:z��*�fv����TtE�Z�P��6�\��c���K��\K!��+���������! ��?[�?���ۻ8�>�ЕG=�+R��MVjuP���F9�S���|�w��yo�����|��&H{� �M�~Zk���Wkێ2G����-��׫�-���+����I���N+�ү�@�4�J�r���^B��ۀ���_Z����}P��E#�05k�+��˰�h	�FV7Ǆe�v���߀gO=�vO����ٮ�!
����:�Z�=	��K�e{(`��SA�'&�����u���'J������-_7���6�w^@WX4Bԡ���z3A������p-K���Yݱ�o�Y�
�tB,�Jw�����fE����SU+��2x���p] ,�1y˜*�9�T��l�T�!/b�2��ƒE֧H:G�� �w����[��M	�l{��Tr�~!(�j��ЬfW��)� ɾ.�S��m��g��fi��Ð|�$�J�]zp��p޲� mY����U����B
�4Ҍ�5����P��Kq���<o!���ãLQv������&�ٞ�8�?�S,��W��Se���;O�7+���v�@zz_��*�������rrD|yj�Ѕ����]�ufԿ���{	�1��E��e5M�F?NI3�܁����u�9
���%�x������\腈TS���q�k�f J��N��H�N���N����1��V�Y����)U�D�V�t�G� h�'�`������U�t8��0�R���E��ӓ1x?��ͤ�٪݊K}������qH�&�knq��))�%�l�� IJ�,�z�Ise�3� Z����0(�.u��U"�b��oǍ	�eT.ϼ�>rb�7��I�8��ָ�㣺v��&��3p��h�Y��(��ڐ�O+��/�0�L��T�\��OKqWy��8&�B�&� ���o+u�4�+"&�z͸��[g?m�m$���8��X/��\�@d��zT5���Y
��a>��#ڋ慒�$�3���#'�&��1��Ύ�����E��Az�[�>����,GQ�Ҩ؉j��g�(6~�5+%	7\N���7��ݚC�b�5�;Ϊ9.�A�i��D����DQ��t���{`�|��<�%lw]D�
9�C�]��=> �䫠�\=�s�Bvlރk��'5�B���c�5\l�����:�d�C���;������6'���g\�{�<���JX���,ɚI��es���ZJo[��B�#��P���fJ�
����A��С�<����^l��h=�}�%7ayQ��h>��#�> p&����ڿ�����:ţ��^�7�]�� �&�f�P�E�۪��	\��m�J�o�p�biRmg���A'U>�*���B�Y�\{)���9�"S�{j���(#M0:�_T�����X��kr:���R;�1^P��E:CnyZs����DEl��&d[x���3q��/��gވs�f��n�oN@[�#c?U�鹹ؐ�v�0��᜸��YBSw�1�I��Ε7.?�^$�dϵ�j	#X?^��%�[��)h�G��"�R�$!�YԗXC��Ԅ%ҫ���nW�x��!I�W��APb�^��J�s�t��A���V|լ���Ch	��C����,�ɤ��d?��d�����#d�	�ԭ3hQK�OP s������tSk{�=~�"As�ߧ�$~�0'1G��"%v$�_���q>�}��H�ҙ�4k�[a�@�x���S7�MRm7z�n�ck��ΰvs|��u�	�����`{���a� Q�x{Z��U���9�QM��F�pe�XM�V�<$�n��1-�=�VV��cs����E���.�US9���Yw��f��磚Q[چ�д��MU�|�11ƿ?���A��Sv�<��͜���t��ej�����	(q���pFi-����Il�r�ƣ�)�L��MsY�Ͼ)t��,���]:�~~�y�B8�{� �8ݛ�~�31ܪ뭶����=���;%�o�Ĵl{?}�dE W%�p��Νl��߁�s��SeG���ZC�u��T'���V��fU��;��-��G�"������EsJs[���EO(�,�Y �ӹ	���@�`�敁���M���uXt�V�g�]=_��=����^ ۿ��O��6p�	i���
,E?P�9�%��%� �����H�e���Y}d]N��RS
�j+��%��|�53��[UtI0��ZR��Q�,���4������Dܑk0
a�~�G�i���|ā�׊׆ ���隬L�v��'��c�������rm��]��:���JA�[W�SWk�9�Q�{NS�P�~���?��E0��@ԢC� 4�i�v�YT[�B�Xa�}JH�^S��USj��Λ݆7���~�c\�y�0.rٜ����3g��\f�!+�K��$�f��B�f ��t��.+�O��Ms4`>�3�U���crD	��n��@o9�$\��`'B��F��z쭒ݓrê o�œ��g��c�V�ŨRWQ8�.�Q�ʍf�3 {�F�)[P��%^c6��
�$��r�Df�l�&h�iÃ�Tt�n�[ �6�� �=�p�9�������?�,�ʹ�9߽_�os��ߞ������j��dX�f��ۨ�m�~������n)7(7���>`�g�%����*)4��^+M��Q���9�"Bg3��I
ِ"�d�c���5i�DX��'ȲP��W��7�:>�\�p� !��/���>cqt�Ў�����o�P��z�g�~8�pd4��v�mU��i���}��ф�.;рv�hΐ��,ފFPqr��d��G�O�{�"���P�`����K@㬬ǲ����䦴R��i�{��5�P1�eJ�g3���f?~�.���#:,�:��a��X���6�;�͌WK
v�a���A�넅ԯ�eex�� i��]�"vւ���7�n�Z\�u���0�*,�g��14M?ɉ�7ޱ�.ѝ0��Cנ`gcO�������Z�m�Kʝr˨ $[Q���R.�>���L�j�7���i+Q�X��;)�C���&���$8�I\R�g�Y��o��>�䟵��SK^�����������ڂ�����?�N�bD�0|���"���}.����eGm׵�mA�1�~ւ�P{�
��6��z-j�w�;.{����'%���ݏ��X�bd�!hS�vu,CqYO6�����T
�6���%x'�u�
��)wH����#��"/�K����}�$��5����\#*=m��G�ON��a�Dh�XeA�߻�1!A7���{_R�"����1�E��l>Ԧm�;x������h�(�4?1�p�����9�M���>�w��H�hY.�%����N�g��^�<W=�r�82%8�;�5���m���<�a�R/��k�YM�[#:��	k�Z�r���B������=Z�iiU�>LU��_cmۼ;�J�o��k�7� l��3q��W�O^�xL$N�_�jQ\f8�T� dO�0����+�t?)�U�]Ȉ�#}~��W'_jM���T�Zf��ӹԋ�k�v:\z��?��C��쩜����h� ZS����M@��ąu�[Hg���_ʗ��)�1,b>x��g�Tm����+fH��Zt������w3p��=gUy�A�<]��q	j9��w���P��̗>S$��$Q$M���jݻB���h>� �
��ׄ�ʞ�+���PP�D�UM�����7��%�5hg��|����.|	��f͋�HB�{�!��/�m�Z���*PK6F�q��@:OU[�C=��g�%+@�X�c�����ār:C	"<�|��W�D1��(�㤼]8�����!���3g*S/�K"��s� � ,h-9)ߗ<�Q4�$�|�
̒�l�F��Lc�3�{͝~x�����,h��#M��Z�g��s�j��<��� җ��P����$�����Ed��y�Im�ĳ�y�������L�Y�����X�b��V��"w)4Nw��Q���C��wZp��/_�&<�pZ�p1o��I�d&�H���xB3��s��d��	x܊o���"A�"�h�k�"�e'�l��s$Y`��c�6З��Z����P���Y����b��xT��A��<J�4O��<����h�j��1(��F��Q�:�����vbƴ7�����W�xG��칤H���1��h/�Z٤�ũ��4��)��e�h�I0%��lFx7LJ��)	� �{�B9Y]3�AQT_�N1V�
C�|���=Wz٢�j�!FA$KA����	���-;���?�Bϣ��wTN�����ȕ�/V�� �� '�97ӛ�-_��F�O\~y犏�㼂:,�|���&�a��S����|B�w��%�Ox�\-��4	�L��d�������(w�D7Ю�BO�tt%��!�Y%��o���r ̛Ĝ��ϖ�(��g@&R��}����)�������ޠY��K�������3�ٞ�l7�9�bZ�s�P-�L�T�t����1��T)�fg�zg�4�v��-�����\S3��Gr�*��A���3[��%�H�xu�!_Oݔ�k�����<��(��FՐ%��=��h�3�.d0�'�ڧVЃ���П�d�{{ۤ�	ҕ1��M+�O&�vg��B��}6�y<a}��0��ح���PK�x��G`�a;U��!+jnn�nӺ�q��J���EQ�M�xR�o!�E�?�nm�l:������sjyX��o�Y���O��=j�F���K����^��^�kBXB��Zqw4Hd�9n�ٔM�+�����������/�^sb�{��cP�v������OX(押�xg��ER�ɟKZ{���׋�s:/�� 
GC5>r]蘽�0�)#��D�6�i3UpJU{\��ƁP�
�Kyζvd��F�3��>E��j�������֜8���k�l	�#���o�iXb�i�W������K���w9��r�d���@�*��"�1����������4�.�V6:��,MFz����Mt-n`柤EAN�i&[@�7�;[�҇�A�^xy�w��F]�jua4���?_V1���X��kX�2g���������4n�j��d8O�G����}�R]���:������E�׈d�LF1�׳NbF�����	Ds>�||N���p����<p�� ����1{9D�1��37v_=1�=�쿦�����N�]�.��o"p�S�~��eէʷZ�h��L���i�� r�Y�MY�1�K�K ������a����q�5���Ǜ/��c��p.�{��G�:��a�A{C`,�96+"*%�_�C{�_�B��j��G"�]����@����:���:�>��o��.����ur묚�C �L�I���
=r�������(��*s����zD
��a�-�Y��=��s�g�ъ[�>#�>0��&�%۪�?�p���ڌ�x��̰�P"��1�dH���É7���B&ȕ�{������D[u.|���*�f�o�+Y��$�c��	�(/B��(I%�?�Ys?\�B�W�]퓈WG�X<�J�н��)�/S��ł'���/[	���?n��#|-ZWc��yj_=�
@`�Ae�A�"�v �xN�et�Z�=�����#�5�n6��L�%"4�v�b��V.�,[
=c���0�!���8+2p���sF��+�cI%CB
�d$ౢ�㔕��DuR�zw^�q{������(����^�qW<� �bF���:An�,V	
mt�QS-�&\J7�8:�$��������S��9��*��GJFL��G찺�{
C/�/AYOZ�t*�qp0�g����Z�#����(�nb)O�zU����BH���E�*頱w.s�4� c�*H� 2C~�Ŕ�ļ�L��b�[fY܁� ��*a����0��P��A�-4.6�e�jQ��t4~l\��
�G��If�{��>z�����C`�rc �Ai��x p�7��|�(��.��ᇌc��=ew��G�A�F�����b\�R�g�����<�Dyd�٦'.�����~�=vY�- v�8_ޚP�߬�.��>E��Y�4�N.��w�V��l��i�5����՛�t��ѝ©�MpnRx�X���;�9c:
R���V}b�(�D�%��~�Sc@�jq���*�T�'!��)qQK�u�c���"a��/�z�QC� ��/�O
�4�1�r �����R.���j�+�p��%-��u��<W�Qs:?c��V�����8bp�ء�M}0�8�+5�"o`�{�a��|z[۾�Oeߡ�+�`��i���lۨ�l@�ϧ�jpJVa���.���|�o!�ǂ�mcA,h{�P������#]��X�0��v�;����XyT|�_�4n�q�Sw3���̈́�{�J4z��R-�!�|�#&v�Kd��dd�aP�����I�[�n�1d��C+����fN��p0)�a�iT���)�G݆�@����xxPR��J��O" ڣ?���{�� �W� �����@�w����'v�#�+�5S����Ѡ�5�)6�z ;\�e���گg8j��\d�?P�N<�E��%�n�6�N�\+H}�_F���Xy��K�A�R�#�[N�BiGKۦϱ�e7��A�t(�5�����Bg���GV�}dY`G���7H�A��!�aaoo��S�j���@��X���-�;�z���!�G�vSqi&�̯�"�9�X?�Z3��ec��S�0e&�v�����v��(�p3�E����z�����[�	�T3�7J��}��g���"�x8��|q���5�9��H�<��B{9U^���WU����Ɲ���tE� ���g�Q3�BiZpZ�W�'��g�/�#͒�]���>���o^�,���W�F�f����잼GLn� �쿁�*�����η�]��aj��$�pf��eԥQ_\Oݿ/]�j�~�o,��ނN+����P9����SZd7��gH!���<�2���Y����ÛO�喃�[�F��<#�"ww�4!��D�s|F���<}R�����'�����مy9���=�L�Qz�! 1a$�;���2��y@�u�|���i8������>���}J̾��Q�s>"
ֺFTÁ׺�T�1�@v�Q��Szb2����ՅB����Wt�|i4)�+�%���8�].��H(]�l���zo�-��u��I|��q���ۋzED�}ya�#�nJ�0�o�ԄUp�wC�}�ak��Gʯ����?�SSK�H��Q��89S�oeG�7YEI�m˘H�Ƞ\�9�t�%�M�F�Ƈ�<�DM�0��\Z�v�R���>�<ʒi�%�a�ޱ���D������>��^����%>z{��`W�g�`���C2����u��VFx՝6/ZB���Q�����a�����}�]G�vj(����z�#��ā&V%�r:����9���iyK������D�xx�I�������+"��rB�
iڪ�)*C��0��C�fy�ֆc��z��1��X�
�-�����t
���u�BsL��y<3=ɱ
N�W���IB��t"���6d�JYS��]�h������H��G�8��5,����tH�>���]����/���q=�mB�_}���u.C�|7 �����z��D�mhX%/���6��&��p?��*9*R�:��B"�nc	����R̖l������A��Q舝�@�!k��W�[�|��6�T�*v��@�'�\��&\qGnz�1+��i99��b��jb���6���Ň��ØEh����$d�����o��;� ��4���ժ��-���0�f)f��2���Ms;l}U���Hm#U��M�BżrLLp�4<n�B�D��!��ᶼ�,��w�X>2u�!0pM���
�����2��ݧ�C�䊢Q������NÆTI��f8�wu&��\N��	�S����\QL���%�H�=�#��B/�&3p82�sv���G�گ� �&z?��.������L����\ED9���h�N�y��X���<T�V0_���L<*)LjK��RԂ��[���Q���1�Ź���	1>+��������b�N����z��Ht-��z>J.�V�(�[ ����+&�%L���]�u�Jk��nk��F�㢶6=��"{� ��H��y*/&�3=���Y�����%���˯l�AFӇ�O�wf|����.roڋ�a�m�3��VA��V��#�/��Z�/���t�y]D�'�5��.�]��Ԭ���V~�f����q²3 ��-T3f4F�"ހ��y�΁��8��!3�L-�x]�D3ޣ����k�����Z��+c�n`����శn0ǒ.Rl)Ѡ%:A�7�,��au��]5!o$�+�!�O���{c����T�p#�5�krT
�$#{�,4�}�A���c<�;	��UE�&ؔA6������� �:t��T��q�Pa�8��*q���u���E�!�Gbh\G���Xҷ�3��v�I��:���d\�i��+��S�	?�;�ӧ�\����{W�p�"�R���8�ΩF�h���ӡ��w*w��ǥ1;($���u�W��V�M��)�Z�Fҙ>"�_�T�i���pY
�ǒ?��;U\�*\>�bsa�v�T~�ǟ�|g��#���uí���/J��!��v�L��bѾ���4TQpdkVXb.�c
v�}]A4ƒ�U4��g���B�Ov'��2�6�(�vZ�T:1Η��ȡ�� ޯ����Uex]e]�hi�
_.��B�SȄ�<�Ćy�2N\�T��'����sv��8$��PrO�~֡�@E�r��w�M��I�j��tW�3@\'��R�j�L���^l�v�r[�|��i�v`�ٲW6��4�^s�9��������_0�<)v�f����(��G=X�,?��%*%�<c7��f��"�o�K�:��9-�1L�O*��s���㟒\<?���(Ĵ/�f�0��WX�,��Cҍ�:�K`�e��nE�Ƈ5��� ��[b����V����;�rq��َbh
��_��[;Yq����K�o�{a�� C��D�#��q��nQ�a<�7�pR]�gRH��"����� �0����5�M�y����׈��T|�Jc�n_����f��
�O���hȤ ��'��r�z��0o�6��ڰ\�8l�iY�������A���	�48ň�
���B��@��^�������������X�w�#҈�����q||���k��� ��L����v_�hL��ȋ=as��Q W�[B
�p�
g��V�Ό�wh<�dҪc�y�gJ��k)�)0=vWh����#��T��o��T�� ����&��Ke�h"�i���9ҵ��A�M��1�z�p�@�����6T������rو�R�h��m���&�n��-��2\���.Y�u���/��B���s��U
Q�7j��ť�o��������Ȋ�����l�W����f�#,D���{-�QdL�aW4<c�j�\�m��f0O��21ܲ�}�q`P�����P���bb':K׵lkO� s�[iW�8����
����LcAU1�<trp��;!}3N��ui[+m"b3�N�E�ϕ�ȔȌ��C"�,s��Jc�4�&�������f��Sz�9���B��gQ���������\�����(Ei�xd	�'�}��qi�[a%{�K�H����ۉN.��P�kR���][�����2�|�&a���T�r�=�ǐ��$�Y ���i!RX��X[i)�+2�wԻ�y~��^�s</F���Q: �O���S�u8,D~�+@H���935� ~a
�يZSB����� /O
�|6��䌪 :ۥQ�V�I�8ZɱK�z{�$8�H��,N�ǟ����j����<&v�+""��XlVݍÑ�?s��[�^4�j���B��ZÔ��.��3�4� SG��iAZMgGN�C���'i!V��%*��_3���[��\Y͝�m@���^ե*o���(��[}��V�� ��$Z�&pԙ�%�[�$qB�+�}�+�^{\��	��B����s�s��q~Y����v�e��	����>�,�����N�3�a�ҷ�(�����12?�6_L���I~�RY����x�_�)>|� ����LIOVQ����|�=���e�0P}	/mZ�ҕ�m����zN��j.ۖ-�&��iX^Q;Q�E��*��zY�v����_:N4�i8����E�+p��zf�;�5��;��Shx$o�׼�a��|t�zu��B�)�g�{O^v򩀟��B�.��A�_�V� �)�`XM�}���_�����4�j���_�#/�-a�2צ��/z�F��7�:_��l�AƵ��Lo��� W���H��Q����JD���Le���,���Z���0�<As�e��}��A��rU�j΁�ry9��j��h�h;�yoWӏ�v�o�5e]C�=��I�d�HC��]�ӵg>�'�8YO�D���X�l[�*ua-�+j�QŹ�&���碟]���-��y�UO�@�C->Bi���閚c������;*?��3t���B\���R���q���ի��f�s�Ktp�cc��M]a��w1]��L]�Yk�4�1��i�
�6�L� �����|3Qxgw�Ϸv��g�����5�BpC���Nd.\�5�v��҄�C9�:��7���k>`��,XM�D�y���ru�>yNKāy�7��sd34%�����)�Fb�*�󓬆�\^!I�w��Y>�47���_���h�3H5�QӢ�GB����-ӠY7�hBz�5�o�$�'�$���*��Ed։ ��O�q�.�����5A�cN�}p�ɚ��?�B�Q��t���lk��#�D��*;T��)m�j�)��ѵ���p�	�<�(e�L���� E,AH*7aĂ4�]�-�F���R !ߩ��X�*��O��y��_(�m�� 6i�����Ģ�%�Ί�}�-�����3;I����8��[�׋@��c�9C&�G"���Sfr☳D�Ԕ,:�Ў��kQ� Q A��~��O 3�����Z�$���[Ǘ5=MƖUc$��R)�2y1}m���,&j�6֦��k�t���-��ӈ»ؗs.e�.�W�y9�Y"E{���~�������m�f���ׁ�"[<��Ns:��2~�������Z�0���])c�v*�:%��٦%�������u��Z����h��̒b#�ڜz��j��������4ɵ� �߾�uw!��>H�)�ӵo#&�Y*~��~�p㥢��89:���lt�"��X���{� M?u���{7VYހ�42ߏ��/}�H]����E��uxk|��,��q%�������D�Z.v�+d˴�w�*r�	U.>�Smw;|�pؘ��14`�`���ì��e
`v萴x����S���ᩢ�-���9�O�Cx?� "����(�E~�kCs$tĻp�U��N�X����U⤭W�Y7��i�B�!N�7DH<�*����ӵ�N
P�jul���=��I�+?�	��+��b]#i&��t��I�-jj����蚍��\5)�.���|���\Bb�0�?��P�G��(�G�b�a
x��+�h�)��H59�e��Hy�H��A�
v�p�u�_�}1:�-���{�G�,wO�-d�����{��Xy�~��ӻ���|����\�e�c��x�RZ��fז&�/hR�#�]T��� U�:(Q���2Ҹ�!����p��9�E-]��� �k��
W�>\D���T��0��T��������d�y��0y3W�1�Ǒb�ŔAo�� Y���Z�od*<����;!��2��B��ˀ��Y�'@��F�Y��7���2�6	���7�޳X韎s����l�gκ"��O>��1�2��(��T�AE����r��*��>�:І	q��	��f�"VgݮJ�t-���̷�
'S�|�=�)���˶��
ٴ� x�g�y`�|V���»ƒʇ��}O<=�A�s9��Q3�n�/�-y��<��Z%��$T����
��@}�d���C�@M<ܣ��;M��HF�9���$Xs�b�����)��y���]�Y_���Qɜ�9f0_H:���s|���ô9�n�S}��B��BZX�.(�8H��|�.��r~�t��t�����3�f�%ʇ�7�"o�Z�
7����m��t��ֵ��^[eԟ%�\~&����HV$�+��L�K"l�
b{]_��;�gb$����F'�\�$Z��q<J"���mV�hl��{���Ȅ���qv
���ۨ�V��"U����%m_8<���_}o�S���M_����B�і�[(��l:&�Bq����О�@���aYl*�0�Ê8V�Od���W5�͛����/�ho�����M1����J�\��9G�sK��mXc�သ�������p+@���-(2<tx[��7�)��e�4��P��Ge:K�m'^�b�� &+|qLߔ�-�����SW��ôf���4hHxk;���U�,�~R��~�$�_����SA��J]�[�d���p�Lh5�����u��L�.�i�t���h�?Օ��o6��*\F��,f�؅��G<?���z��.�נX�9��U�O�=! ��D�����G�7�M�Bٓ&T�@za�H��ɟN
�mHԲ��S�w���#6�څWG����N�]��w��t1l��¼�8,GW)ކU����g��F6���֠T)��atd�zf\?�2���y���r����䟀����O޿��rš�f��Uz�i~zk`�$;�����;1[(�_�7�f�"���P���uz��Q@X�&���ɲ���|�*�-[d���
	n�hc�3Ɏ�u�v�9h}��>�`N���*fuR�8�熿�g�*c�PǺ����}�JA�Da�heE��R=�E8J44�mLpƬVG֫Ep�yowV��ڥO�6�B�ߙ�ś4����Ua��(:��²���}�?��d"�E�"�H��v�g1�Qs�ъ���9{�����Ab��}���(�sW�T}t|'Agt���i��$A��	d5���X?qbVI�V{�`�n���#\�G��R���3T�]A�򵕛��F[�q�C�� 9��f�{�{M��l� xH�.	F%�rD��y{�JTBs��볕����yf/�(�=�2�J�Cy��F�{�o�R�X��e���L�I�,�N��j��&�s!��ˡ҆���S��`�p}���!c�/���ZՁ���Q��W޵>�kg	�X��;5�F�oC���ㅫx�O��x_,	b���M�"v�¹�B�sv��J� MY�	�A>�D�䱀`8bz%�����y|Ya[��fI=��ꥉ��'�*u0�H��yV��Z���S���2�yj��U��u����xC��y�u��Qa^[�=� �5Cz}�gm�Wd�[4�[(F�rMbl�����As�Ѧ������oCG����kF�E,��y�ɖ*6 ���z�.B�����(�f+[�s4%�W.\�}}�g��
Qg��|�2k��g�N���[PH!�5!s(�Y\G�,ۚ��Ӱ���v�ɂ�?�X%fy���E���{�GSȠ�7�g��B�|�.�v#�ze�v�ߔClf���d��C�%X�$F;��k�48"��*��P�_��1W%�x��!�������mI��ف:G�;��")�[�5f���
=W��s���2�\�C�Ӈ��>z�#�D<��:^Y\����	���h���>
*!�6YE�Ḟ�'QA��@,CN�JC��ݓk�i�K8��E8��F�J��	D�_�k0~0r]v-K��$x�_����%(�W �k��$��k�,�֎�؍�?�[��R������Q��fFz���5�aZ /~�у�6��ȠI/�G=�ҥ��k�+���+ M{�a�d/�{���k�?��.�2����6����q��?@5��QF4��r��� ��Cm>n��6r<*����=��)�+��ՍĘ���4}��6�nX�q��>+^�'����/�i;N���#~�p�&v�#,��ރ+e���~��A��R�"zHEjb%�h�r���R5G�|F T���ɒ�����̫̽b�Ӭ��৸@Dj�L���8��]���g z ]�����϶d8��p��Ok�է��� ��_�kN�0������̇>����(�r
|�3���BV<���>�5>%��/ܜ�|6*5N�)�Z�e�����k�g�",��0B�{b`���6�� A�ciϞ�0	r�����`�/�[�?�_����I��(�g����XաU%�P�����)�Q�P�"��<2�D��� �.�$]�^mŰ%�t��73�3�Q����"q��_����h|���}- 9@j��Wqx�q���y-�K��W����:)-����=Ml�F��z�5 |]5�U�g���*+�^�~*�D���7�q׮eؘL�2t$�N$Xݫ��@E%�w]�G�|�p��yd���F&�uxI�V��좻�b�����i
?D9�A$�eڼB��sx^i}�&I�se�(�T5��J4�EA?T��:�V�n:(�y��l��D���4]N�3�N�9^�z���n?���[���&2�N��rY9v���#��}M�igʷ��J�Zu��J�]Z�vh!��G��m4Tb\�~vN�W�^W�f��8h_�������^[ eڹ1�^�j�3���
K�W��+�u���/}�����;7c�����%�D`�����o��Nd4��nY�^�Z�]�F�es��A~:�!����9[gw��D�@2��+W�����:��%c`��%��ƆFl]P�'��}�/����0����bfW�:�v?�0���X"�����FL����(����&2	�/��u�e��?���<	�!����NM|�su���1t�oAiH�o���}(�mx���_�uVǻR;,7e�C]?�#�E��__.�l�>
!;[�?��3�v�hx�vI�Y��>
�k�'wݦ����9��ڳ���y3o.W�>p�w����>̭r�1ak���fh='�]����çCJ���"lH��vrq�����9�GS��#|@�#F���Yƾ�
+���e���f��y�a�p$��]�襣ɣVTbr��IT2G4=C�CU:���iĄ�U����Y�ռ��Q��ҟy4=J��j�����g V�����b�7�Z��ƾ0�i�# ��LL��i�S1�[ (��)5W�3��Ud��#�I�t�Px� �]+� .��g������V��&����;��Q0x�������tnW�m�7�hl@����7p�S�6�*�B��n�� '���^t�C ]�d��H�c�r��~�V�r:�^�[�?E��i��|�o���-9����1�FNUk����o?:{ZV�?0��Lݚ`�z�S��5;��^t=�63c�=uFi�og�G���O}[�-No��߰#��.��*_��v+9����p�/�����K{䖺`��y����~�/�bK}�g��";�wN= �Z�Z!w�&EGT�Ira�X8\�j�h�7!`pxŮ��\a_ӣͨ�B�3E����{�!�4?P�Տ�	��<��٪��n�X�ײkrE�K	g��Ϙ�L�0Z�_8f��mj>۬ܬ�&Y;�����7��R>"&'z0�]�`������V�S��ͅ�¹�1�J��Kh0O�A�,����ԯ�.� �9E�A�AT,��x!��'��۝�A&��"}tq{o��1�c�
TՆ�y�ж�Li�����;���܈��6���U�C���'�j�X
�.0�U�"҃yT������g�U��1�i�=ҪdU��1��Nn�ɔ.%l�����,F���}x��q��InR�[�+Ⱦ�fhv����Q�_{��I�Xp8hd�
���)��n0xӨ�_)��V݋�@'p��:5R7�XQmm�X�.�J��rF���h�vӫt�axp�(�FeN���$���S��� ��E<z�rlF^2�w
3�+�1�E��lD=f~��(f�JqL��`��t�E��z��#����A�C?ł��+���i�-`$��9W
jE�⯉"8���U2݉��A���䬐�l8�w�2��Vx�g������?=.�؇�!r)�)�WI�_�ݸ�r�]mO@e5F��衱^I���J��ԣ��J8�dz8w"cp�g�2� ����"O9[~�$��O��}�Rَ��0��{���ׅ�UY"ǌQ�|1AMN:x�K4r�yY'��q5�Oqx6y�Ѭ�L�^�u�TȐ&
�<��X _��I��oRإ�8�X�
m<cz��M�7���	cZ�Ҭ����#n��vv �d5Gx�"�NɚF�����3�sG:y��L�_-����e���`t�i��?NL�j��3�Fq:и�>)�uHFk�����u臰������)�� ���z[{ϾX%F��^��c�|�E\֊���Y��?B(�4�d��-��n��O!����Ɠ���^�h�3��,x/$������%�T�5V M��y����7cn�9�n�����s�51�hS��.$�Iqٗ��j\�+��z]�F5�"t�mn�Z S�=��1b�£Y]R�z�r��*�cU��j��+���ۖ��<���/�|W�;,X�/� �(�c���y������} H��u4<,J �;u�+�+e��P�6�J9�7�Ky<���g�)��~
h�h뭫+Bϳ�1�LN�������T�E>�9TV:��x+�k�f�*�h5$���uf3��k��[�n&XX�01�U��a�_��X�"%{W=VGB\"'2�"��'?U��}Unsq����2��vYnS��R*m��F"�
��۶:>��#(]?�t�VG����ĥ!6:x����fQ <bH��� ��b�t�d���� �|}t�b�MzW�#�c}��/���� `�����嘯��[u]˸����'wwi�l��f����+>��VIC�v�u�%���#�R���!��C���7h/��`��2�޺˖��J�-�Ol�^yF�|B��5r���T+��/ֻL���7w�\�0�3%p�9�g!��	��,�x훋_ݺ���m�Ki����'88"��Kcf���ţ�/K�q��u��p�������O�f3 ��@q	:�� ,��Ժ��㗹/����㴭�_=EK�^S�a$Y�e�ꛈ͹k�|�唽H���*��7r�G��2R�I��킗$h�8v��35���a ���ޭ$ݹ���a.	��>P����&CsPA��\�!�{���<���eW�!:�<��y}2�y��F�//)�����7�W���i�EM�]�+�CnQ�x�pa�7̆����.w)l�d�U�M��2���v��n'r������h��g�k9�,v�LCA'������ҍIYmϏ�8(�g9�Ah��!��R�L��魳��ST$��:��������%8	��
/S��,���3��G[S����<�ea5��G��LB!1g�W).�;�{��׏�^4G�3hUķz�R! � �ܲ��?DF���rA8;R�c���
j��qʜʄT��FBD�gɄ������޻7H����?���qO4���a�lܼ�I#'D��v|<@(u�U�wȻf+#�M6B�2/�	t/Z��r�G� ���1����A�п;��H������yD���gN�D��6���P�9QR}d�ո��#I;�b��/�3�L�X�*4NbԭN�MI����(cy;��u=�FR�����n��q&�m�t�.o2h#[5?-k��w�'�U���[�.H�0DHTw�?N����}7�]��8�;:8�au���m?Q�8�k������>�|�����,!R���yX���LZ^�/1�ۧ�Ug5?�ΐy�`�ˇ��<�)OΝU�y��J�iU��tI�̉��N��6��gN o8��H��2�C�o/�BAn�pMF1c�L�����%�o8��b��4H#�e5_�R ��0%N�}�M��(,�q:.�)���vt�����h�Y�o]�B��%�K����ET���_W��
`u�	�Y��}�����v��sH�������<��)�eC��xi�x�_�tPi�Co;OY%i��9�q���d�����g��C�W�\/�$�3���s9i�s,W�B�#4׸��ٝ6q#7���i��O�n9�[��@IKO�n��d#!?l'��9�U��2/ͨ�\�HbD�^�g�/�k:�xNt�iF�|fI �6�<VRO'�޹�'UԠ��z��Ďg{�����o�D|�V���m�k.��h��0X
�Q�9�� ����!�a���8}o��we/��̅ʳ�B;�,��8.���c!��g�������4�OJ0na�I�&x����!^�Y=�o���op������E3�Xd���>˟�s2�i��i^��yޟ�|�uw�8���H�� ��_rjQr���W�ސNb����eI�5:�^.��'&ľ@фI�0�+��.�,q���=j/��r�ߤn	�׍?p�l0�s�%s9:^_����<N�:(:v�-{gU}�H�
�	E�E-����`"����"+2�� ;����{�ۈy��eY`�[�'ϝ�+�o� ki��%-e=�Q�8�$��1�|0��v�4���(��$?cQ�,c��L�n�3ʫ�,4�Xp��^J����[H�k����v9>��E_))�8ϩ������WlP�O�q" �?�qaYxVtD�Y:�m�W+�G�]����,��aF�K��v�M ����>r�2�w� �~��'X������	D�=�o�N�\�j�3$=%�@�,��;��*�ʑ�צ�z6�C6w�z�ظ:RS��Mc �"��̖�K�g�!�]�B�,�����<��큻غ�� k	���qk`Q��nzV0�o˫���=<�1�vV��ǖ]�G���F%{����@S���i�?���(��k�i�\V���x���R >g��M� �A�����?)���8Հ>34��87T|��6�E2�OKi-~���4��x~����	��7�B�
9=�W�OH2X�JG�%�򱯼l��	�E��h����� ;|`g�U�g�\��T:���m���9#sZ�9�{.q���!����HP��Y��U#�h�Eb�eIv3�8��C�G(��@w��gItV����9��5�4$���A#7JI��r��*5�`˛1����Nh�"�ʯ"5�_�V�p� �z�iy�YҌ��c�"�NS�yPwgZ"�.��q�8�}cp��ϲ��w���|���4ꑀ�=-�JB ���7���S3#ë�v���rs���s�_���(W�������-*��ߑ�d��I��S+�	[̛>�X��`~h�!�l}�j��3�PD/�.M`?�Z¤��13��T8����ke��f���-#5��a`2�;��0*��7����W��Q=�Y�Co��)�����$��8<?��Mv�2f4֨qT�g����Y����=JB*���Ҹ��$ӣ�p��pm�p�wH�U��Q^����$��]���Z�O���5�LR]�4-���J�qה��J�S�f��QU,B�2��\��/Y�X-�x�m�,�}�`�ac�9�����E��6�Uo�2D��!��w/�s���/�F #� �v�0�����$8B����>��F9��ɗz��#D[��Ŵl�./E�Mh��2�� �u�{���ՠ��70��$T�$���{F�ױ��.a.M$!?u?/f�1��!�s(�hy6�nq�xA)����?�+�|�!d	�?ū��W�#0�ۘ�^D�)Z�x���cX��ϚIm$8T�0�	Q�� J�EE5]W��jwA�rm������g�F�M[�9wA����X��5��
c���G�<��Y0��E����w1� �Uo/�s�$Aϟ���06�ϳ��ad��p�!�G,F�[���7������r�i%�������R���^��YAZ5��j:�6��w���jA� M�و��Z��l�q5�K��<9 i`%6}2��v~U/���)�3�n!�!��V����ͻYZzATr�j2B�)��ou�ѺbnZl^�:�hOH����u��u�kH��1?�R[&1��v3~��"������C��@7Pw�k��/p���E�*_���ZL�0w�S��ҷ�x�_Հs����pP��Bw��3�����6�KD|��dFD�q�Z죍v;7aN��j�l�`�~��>�e։���dWH~m�9?Զ�CA��9f�����S�Z�T�<w��8�Ʌ�mƬ��N��g1J"{۱Z>�؋^kj2�k׬Y��E��D���Qz�`�b̎�S(ۻs!b�q�j;]I��r¨�*Vk
�â��ɂ�����]���h�{�nK�7�N����/�9�8�<�(�N���5��Qˈ�x����KI��`�ı�]+h��,�v��'��A��A����{;u9ad�5����#H�3.0P���u$+����e��y@=�����oT\���o%9s���r����3q���/pvK���L 9�ڮ۩e���X��qV�A�τ�v�����ɔ-��P)Ûͅ������!O_��<�\�QQ�� �����LY��y`�첊�̦�8��E#����l!��ꄾ�<M��ƴ���}�Z���м�/K��o�>[�xzJ1��u{�rWjdz��6��^wI�U�����t���`�P��t� |�o>�����E^�dʊ\�0Kv3qHxx����u�@��7��~�A	*���iXܞ�A��u-|�������I�
8�\<WA��}K�A$��.����c�Q;SqL��]#��
����f1�	�B�;�D����qe*����� 3'���eD�uZqE�Y
'����&3�Ȟ�G h4ò�k�:D�l����������N%К�Y�#�6��ʈ �;��\�K=�/$�������fNa� �L��0g��2x�6mm��Ι�.>��BpQ���b�x�jI2[�V%zpڞ* ""�P��*��j)�=�k���$0����G��Ĕ �t�[�(�/���P��C�^̕����4�`�8�U�_م�S�7�[��,l�h�%�|�1ɻ����<y|�ĺL򋃫C]*Q�����F��pr妈K�d� �r93��P&[����@���m��E�jX��,���ϴ�����&?�H(�HK�l�OA���g73�+��XojW{$���nœ�l���9s�yחY��´�LE��5/_���e"W�u��)�$<����`��ӎ㄁υ����g�Z�:J>���P��j���!���^���Ɗ�r]qj\b��ǅf��	�^��z���(;0�g�:�+ӳnQN�r ���[��*�ZrzԆ����'�S#����	��F�����[����-|���]�%	Yk�����;HO�Ky8�2sy�⑩ߓ�LW����@�mdwh֙�hxG�Vr֦m�ǩ�f�A  ӄ�
l~���`��4=����}�]��ts���pc;pΫ��,V�Y��\o2��}��
�h���9� y���(ε��ԥ[���M�u�if�c	�����w�H�@0�<��5��'�����w&b�=��JN[51����{��
b�������GO��/#���I|(H�}y��4r�X3�L�!*�R���~��b��c��Ja�)=�����O�#&�T�:�3z�Aow���,�ܡyؾNL+����2���L�L�\C� �U��]K�~p��$�C`!�zO��}](p*�|ˆ_�EE�0�R�BT+�'{)T�U�Ri���~�b{,�[�%�G�9<+��H�&�B�+ꮕ,��s������/�ŜS���8��M%+�]�J��X�&c�g&U-U�U�:5� ����:~}���]�(�b=B��Ui�@z�mF��Cru��Ϗ�	m�#c�	{�������i����T,�Fp�=pG_z���I��z&5�n�7X ��P{(�zY��x\D���ʯ㻏�?A���(X���t��r;>�kX�u(c���\ ?I9&<�3@�7��fj�b�\�'�����-r���k��䂚�}��:�������$	����I(���N�3���h^�2-�fQ{~�jáɊ֤��+�2�A����3����B�,v����eO۳u�dDB�����K������#]�~���D����?�;�
M���^�s�DvR(mJh�`m��|�6�o�xI�G�=Y�k��'O٣o��6��*4�}F��jI�������bDM��v�T�5�ъ��|�kaw�wyt���dd��T&���5����eU���1�H*�؀ؐ�Gx�����b!^�ぐ����#��c\FS�"���� ���߃c��n�vl���28�����`(��0�j��De������X�L���\c�ܥS9���C�����cK&Q�BY��}��/Q�F)_��b�]��?�[�e�܈�[�V���g�tOk���s�*~�
km�X�۞�<��ß.�ؒT!�|b�M�H}`l��V/@�>@j�#H�$@�>D�i>��FlK���#R��>+�Y�i��Lm�����H�1�p��+d*@:�����y��%����������`h�9��N�Z!��6		� )�W�F���8}}�9���0.*i��Ѫz��(���p|9L�Bk�F��$'=��"i5}��Z |/�J(ň�'�f&,SN�Q�~7B����Q=�D�_Xq7�|x�k��,!��� �Q�d<T)�VH/�4��ˮ�\���X�h<��M�7����&#�Ɇ��錼�9}������{2���M��R����&Ɔ��߲�Ͽ�)�}3-i�#,l�{F��A*6Ͻ>(�-��϶��E5f_��A\�Fi�IsJ=g��^�ք�F�Q�-KkH���0ٵ�z���]�ό��m�gz��ЧpeC���" �o�d¼�a>�y�87%�( �Js`,O��j,yc��3F��օD4q��kb�5�bw�3���2��~�ap�xo� �J�>����:"��>������am�"+���l
�]��ա�D����L]����cW�\��4�w�e�g�������q8�CZ,_6F��W��Ϙa|
J`'2�dXjo,m�3���]�JtLjR|-�؛�%�0��k4��<�,��;VL�;�9�`������HȽ�_�b�aե���˃���ڹ`t��"���^dU��~���������;F���G���9�у3lC)��.��ޙ���ҵIi�%�O�ZZ���V��~�F3�)�m�=g5���G!W/U�XM0�M�g����k� �+�1�)�g@^���P�.�����ztK��2�G��Sy�O*��P٨?0^��Cg�'=w#�;Z��AM�Gc`�:���}�U �
Di	�mȗ+c{��U��qiO�J��:�u������0�����L������į���������bH������?�@-K�D�`�o"��B�KW���C�>����&3�D�yTEy�sa�����?ϭ�4�Ab�5і���|�p�����1�h������)2*��,ӵ�xDV��]� ۬k+ F{f�6h>\��4۾���<���b�T��Fb���
.wG����"!(4!�� :��bN�.m���}p*75������G?(BD���K����8r��|���J���/a��M6�"�LuY֘�kX=E�CAk�b�;�>�)6;^���,��<���\j�E\��K�)|D��Ӥ����[�d-���jx3m�=����$�8.n��<ȺB�m]M
�E��RRe���I�^$�k&���HL���)�C�Ad��>�����cV�n�	����Htc�S�Ql&��D'�����vv���lo�H�3��a�N����-��E�pIO��GZɷ��̣�G�~��[K*ꡝfS�U�wR�9�&L��6~#�0q���&�}n0��^�[%�I-6B�Y��o�
���>.���?G��Y��`HÃ�Yh�(ۺ��,h@1'7�֎�����yaz��� T�Pn��vq�L�+�в��6��i�EZ'�8{��C�k�����:���%�qs�_ȑT�����
D!��ђ��c�4��=��v]jÈ�>2��w��F�5�"߽����s�y��ZG<�C/ �����XL�e��F��U�w��uW�Ŷ���p>�&!��M2,�B}��Y�u��|���
 �o�w5�����O=��˭u(�<�8��q�l�[wfi���y��(eݢ�"�͡����$��b��R�l���f�Ŗ9B��A�:'�F4߮�C�\3��
�>����6�C�[Nx�k��6̼�����8q�&!u��Gh��=?�� �\T"mXe<������i������I�2 P�O@�cL��������S!�q"��~{�{�m?�,��Z)|x��_*��c���h�������31�P�e�M�AM��Jx�Z���y�9�O?��G�G�0*k��
#�T��J;SSe�3���R��x�x�`~q��zk�I�@��7�d�&�uaA����E��[�ۈ�<��"�a0@�5
|�^���MBJ6sB��{wgU�����E Orڂ�ґ�l�q�wpr��gV%}��8h�����Ҵ&��dO�E��nD�ɖ>�H�i���	I������V� �q߼B�&���'[e�\\w�8��*�!zPv��?���&���`��$�*B"�W��'���ǃ���)e&T��_[|Aԍ�4�YO���tia��U��lu�!І�Z�����[�+��� ae�+��7}���6��kE�yt�6f�hZ+�&�A�E� �RX2�5�;�`��=����?$����'�4J�R�����s_MR���z�ߖ���I�����1]�t�Ҟ&م]��zd߲S��p.��=����ia�}��a�1<[:����^ƽ�+Rn,Á�O���E�����5��
���U��"�K��Us��ҁ�hn>�������΋(�+:�p��݀rkO���4�j+U���M�I8�1���GpR���BE�J]c�(�f ���n)���[����+������vn�l���C<<�,5��~�{jօ�����Ί,�C0�]ԟ�k�T����a��.��Va(>����g�XS��������&�k`�l̕6�Xu �}��J�<�x�M��>ӹ�q��>�x[�j5��Y�׮Z9��L���r߱��c�1/�Je�U���(<��J����ȅYS��`Tg��B�R*���),�r�uQgE���ҵֶ>��h�c���T�rb�=|X�}�@�#�ǿ��oeƥK����e,�<��-��!M�)�m���F�6������ĺ-�-����:A�+�N���9g���̼!HW�8�����҇
�`�_:5�v��P�u[ĉ�M!i;�ƾ.j�-��3e:���4Lu)�\TqJ�/�{;%Rݫ���H�wcY������jѤ
����V�IP�Ђ�h��>�Ϩ��L�=Q�R\�F��8'd�i�&�߭p��&ʱ�l>��\I��d���e��a�q��@�tV�>7����:N�۰֍���1 3^ /�H��g� 	�E�e�� ��)%I�k�	��"��X��s�T�LE{���R��1/�ĭ@3W��x^<��Q��P~���,̲�����l/��XS�-�9>�ܲ�̔��bױ�1�'t�t�4�p\sm��L��Qcg"�6�����Lt/�H&��-�}h��k9���T���W�Қ�F��h�p$N��܀��Îv��	8/���"
��n Fu�}ST�����gm���'�4fÞ��(�y���栽c�����̱��F�'�&S���&����ª�@X8���V+��_T�K�w��R�!�PFQ�M�
�D�qS�J�RNR���Q�^�t.�!�U��i)�ϔȕC��K[+Ќ҈��������"�`N��1y�wif�E�4���\� g{�cC[����Sy%&��6I
�+n�{^��;@y�A��vrM�ȡe��̕�#z�Ⱥ�'��ȉEYy�&k����n�~���'�b�/i?��N|��Q.�	^���w�#ZM]g�������^Rg�+�\,����P�I���Ev�1< ��θUU�YMW��̷3w�T��v{\�_r�r0:��B����r�%��]�<��1��v�Ȳ@���X��)l���{�y����I��D����Iu�hp�G�I��P;��o?�:�
�n׺g�i��ٽ��S�y?�F��a��U*~,�í_���8���/�;W
l�ϊ*C�����#��C�T�jF]*d���f$���L|��֭`�Tb��D]U���9�7�����i�]ϖQ  �L�v
��@��ntOO����%�����{Q@$���ry��k�/ z���9y	= m\�о�vo2a�9�Yn�n~�X=Hg~V�];U�H9����D@Bo�e�Q� V�9��P֘'�Xe��/��{D� �U��B\�D�B�w�f(��uj�U��ϕ�����8rʌ@D�K���5������W��wl���Nb�"�g[;S59�ˑ�}�2�5����G�}\}|�uo�YR�q|ܳ��Śo SOޕ�it�@�[ �M��4�c▟��NMr('�'Tk	�P���ǘo����9�[`�0[C��P&1!;�]3f?�\*�u�w1\��C�Z;C��'��#�*z_
��_K����1�|,
z^�V,
ʒqXK�E�,��1�32f��Q�D7��08Oo=��IZB㉮��g)�R+�>S�+��[2k�c��=.��P9d�B��7��Q�*����v�_���[<�a%-��hԬ"����b�AG��Ɔ�z��įuL�͸U��[�B蚛��8�*���}@�c/�z��S}����h~�r��2 	��f�(K���&��Y�����ks�i�	I��:W��;k1��'@
�w�R�}c��߯�C�������!�A[<�%ص��s�`�.��͑*��Q�t�k��� g��D}�\�#�yPL�Qw[�2�d f��7��� q�%L%���4󮤎�Ȩ�e]G�~wd�V����#*s)j�4ӳ�k!�'�m�6a��$0�rv��twWw��8�5��V���P�������c���ʃ�� 2�����5�~S��U�AJz��GY{�p���n����f�H���&��r�ӓ�J�۸a!�> �n�YQD�3U�ӳ��5YJejҋ.�vE�����T�I��	$�#Olt�s$��j�����	�v���	��/��t�m��؇.`"J VV/��>�iZ���	b�F�M#4�#-f��
�(�cv��*pN
g�W���mD�w�/��ǣ�SP�bD��84�����;��fSJU��G��jc.�W5^��h������k������Zdz��fI�i�$�ӯ'���m��f�����xš[�=��H��ʅ�����������9Sto�1Ѵ+��Q�9��}�xy�:�ǆov����C`�sU=G �����:�����@%X�O
����u$<�
p���OA<��q|��eX����ϕT���b� <�c�@�E{Ƶ�<�мG�5c��dyK���yI�$�<k�5(���6��E�ȳ�q�a�XL��@G3�v�)��~=xm��	�(�m���ƥ�{�8� q`$ ���[N��[^O�� �R�	�(1Y�V6�XE/#x�?�=TaT���<�B/�\�����k9lQ[������'KX����#�;$^���`SBqt�H8�ZU�I���T���)b��J�{�����?-�{�@�~½)��Q�:R�zG�Ƿ���M�>�,{^l�>M2��ڲfaZ?�WZ�>�U��rMMd��m�qp�����zZl�Y'���Q�zg�
avh����2"م�!�z��ui=�������e����Y~�UBuY���X�����a�$H*�5��y�C��)��¤�1з��0&�)�_�Oj�I��cvks�]�dxI�!���";�U'�Y��.���|!������
�m���ҦpG�cpp�l�c1ޅاS�i
��_��P�z$%͗�4�xi����#�b����C$	���L$���ۨO�JfQ���%����<���(t0�
4�r�㣼P����e�	�č@y�\"�>����%�(��3��4�j�T���(ݭ�QU���z���Y���b0.��7њ�s��pl3r߶m����̨�	�}?'�$��� QX����D�SZ=��̫wb�l�������df6�t��Z�Ōw%�]��*G��U#@�4N�8�H�|@�)��1Q�W�,�u�]�(�Ҳ͝�u:A�����G6��|HhP��L����XK����"���7��!+[�6#����Jjٗ��'�m+�փ>8�<����!�v�fd�+���}�a=$ ��2v����Hk�7��^X�����f۪��1P�����F��V�h��_���gs]�`��,;۰{꟬�9���S����a���E�z����	�)�LT_��99k˕�����}�K�eN�Z��20��v����.�H~Y�YWHh�ď����i�Z��8v; ��/h��x8�Z��,��-���s�^S	I���׹%����.7���9!K�9��8�X�����)A4X�,lk"7�"tN�@�n��C���c��o�حK �_�Y�����H:.D���b�s���z$���6<ʐu�W��ô �x�ʒ �.W�#�̤R��S����'���݋a+�/���ڭZƱ#�.x�����Je����������rd 0�SG�1"�Bj��hR\J:$���yf�s%�	Mv�y�rN8���� 85LJ$1����:���T�eŶ-�z2�"���B�N�����;��N�lv��u ��e|X�+a��+v�'y�ݷ�f�e��Ȝ{�6���(h��|��ly�Q��Ȯ��ل���Ԃqr�*O_�n4��)�4:i[ޙo��;����/�B85�X*�_��Җ���i����ϰjr�����DP��:���!�g��z[O{*7��9�oṠ�o:%j�qV'�qN���L��+���=X��Я�{;Ɲ��K�Xܐ�ؙܾ~���c���5!��[�_b��q�N���,��4A���VY7�:.�$��Ci�\��C� Ρ':��M��Ma h�i��b7K%�����a7������lE;�4���*�U�MV��������1������T�7V՚+ۙ���p��s@�ag��ܤnu��b촄����0���1��,��Z*9��]��JϺ�Č,`(e�n��I^�ҾBA|P���)�F�@�}��D�q�|�ThO'ϰ�x�';H�����S�J��^eo�\l\���'�R$���K@ � `2b��P�Etb)��� ��l���@|��j����8�&���m�?H}�U=��������(/�5 ]o�G�R��qgD����B{L���x��F�^Piqչe�ݠ�GJ���:��A7��yv����y��Уr�L�,"�����3�1�[�Jn&Dkm���n)Ӄ$n��4�#\�,�VN*{��Ir�C���+��<�)!_1��,�Y����ur7����� F��Dw��"/@�=��
?TY�e[��B�};k�O�C���������ɦ:]�U,�_$E��DF��ɂ�%��;�V��o�2kWzi,_%b���lh,H��l�t�~R�ɷ��{� �Z�_�hq"^�ftyB�eUè\.F�:����D#�C��1&N�9�H�<���ݕD�V�E#^�_u�n�ވ#����\}�]7	k��p�6�]F��W�X�,�ZB=��_�G&k��~؏�� Vn�ϻ��b�j.�۪���/�}z����Yj�6���"F���qѯV
�?c�]�^5|ًI+8��M�PŦ%v�"}%f�)�1������W�v�)�!~�W�vik��k���r�=���K����) c�U�U)m�+A��H�����L�G@>���p��I��2��v���ɚt;�C@���m�u�'�Ϥ�1��wCF�����y.�� 1�}l�c΅�x�@�z%�|,a�u<V��_�4(aO^�!� x_F��H��1��u�op�x��QE�Zd�U��bjw��W`���s��Dh@��V�+���Z�V�n����<��?b+�bw _��A�_��׆��.a5~A��~i:	��.0�:�����a�k����<ɔ���qjm��{ńXY �=r5!2�9[D«��O�PuU�1��*i��{������4~��8p�`0t�K��d�Q��va��#顜���'�����/�VP@�>b�b�~-h}v-	��껺��ݭ.�a��'`I e�N�����i6� �����{���@�vŅ�"(�.7[�ԍ���u��щ,���.qa���,S	�{<=����pd�R1�_C��v�ts��������C���<��b8�K:?P�i�Q�5�_�P<�tUN���!�<�@橪�����G?���^���G��6���b�W�������[Ϯ����%ig��H���y��L�y���u�҂ΗHﱄV����������N�Z���cQ��9�J����9ǚ�	t۰���x���X4�K�Ȩ.�ƙ�,8�Q���@�����L|*(�8/�5��=�{}�j�u�g=�J*j��ι��Hkд��gpn,~�A!�E]k8��Ɇ�>ͳ�N���1��W;�y�̠��g�����U��R�D������E���K�:�Ux��Nb��I� oU�e�b~i��%��|@Kh�Y���R�f�"
]C�,W�_�NL�2f,�>�^�_�����{�~���瞴�j5���ivC�6 vk=0S�HXrW3&��Ϳ���Ї�ܕ:��S�Y�
I5c#\�G㡂��-����k�_����?���md�҆�ɻ[�Vi�&m��$S�9��h�V/ż-%y�#���0]�D+�T�7��M<=�ٖ�@�}&�@bE7[���acc�+���I��R2�~:d��T�-���]�v1�U��#���0>��?��)31�VM�d�k��t]�U�H&��$�2é��Y�G�{���D��#w�e`]#t���P�h.��e&�+��"[@�w���˙������z���C�>�{�v����d��g�&�+V ��%����i�@O/��F�C�Ց9EPG��$��z+�r���O�1�4:S���(��w-j��뿐r������2���³��H�
+(��Jm��J�;��-K4�D|g�����{�߰�xi-�惂[o�b��KO�;���qW�����E�~��P�7RBO[qC�/f��l%Oϥ�_'s��|i��A��k��`M0�2q�"L�e��b{���n�ʵd��|��6�	��d�K���|��@%�c�Q��� ��.p� z��Z%G�cX�4O�૰>�s�F�#"xxY��%|@�m<ږ �hh�`�L���[�!���S���{�h�l���Um9�L7�%N q����V�+����b��H�^��(B�+m�����*_W�G�mUQp�
��ў�[)�B'A� 9y"���Z��
�4ah�x!k�����ԕ�4M=�����,��\��22꒑�s��I^��؜��k�jg�ҷ(��,��H��=��f���d��CN�cD�9�����܄d�< _O�B�wU�U�bwa�xւ`����bT=z(G�Piқ���"i���V,�KFg��\�+��8m�	>��cQ�����h�f�@���#�?^y���|��*.��n$�`��AN�'D�s|���1\�浓�mYq�mz��\O+qy2l����LضM�r95�vX�+\{��@(�ߺ�KYc���`�P���P�H��i��V�6�Z�����7y�P��� ���4��P0v|�5	�1��-o����F�wI�8�?�6��/S$Y�������f�z�����W*K�A`�������fn�j��YvJB�:x�ig|^�yo��$WCr�b�	���8?3�y�N�j��0��.Og�±��>� �>]�X"�Һ��Z�V_0�jB�>�f�p�f�����{)��M����%���$N
͔�ƨ���G? :XYѓv9�'>\�z�ǣ@�{���ͪ��lPG�1�F�00��c0>ʴ^�y�w�i.�}��?Y���i�Y�9x��>�S�\*_�`�G/�w�r�]����g7�������([[�@�'M�����h��E��c��oA�mC~�XQ.�GzW�3*RH�6�� ��Oa�G��;���N	��� �����@��Y�>���\庪?��Ĩ׌�>����nP�� 9�$X����tL���]UkM�-a�b�9��I�S�#���!Ǧ)q��?���ǅ�p$�yP���:7�����x��P"g2Eu$���/��w�K������|P��[�@5��h�jTR�ug���$��N7�9�:�N��*i��;V5Ƥa�0z+���|L�?$s[$7k�ER��ͦ�݅y�(}{f�U����ْ�`�]�毶i�6:lz���%���N|5Cv�)B���Q�ɟ�g1)�=�"�1w���$��Ym�_1~��F��򛐭������_�S��G����d�S�e@W@R���]-d�z�&P{�j�	dGd�}tfT��V���@q)S�5��Ɍ13���Kvr��"o`��[e��n�7w��kY��������0�.��6���U}��%U�Y3�L�ݷ���;+�� +݂���3W��EUm c��S������s9W��Q3��;�Sn��j��+|�ܪgu1��#����bxMjq���Q����G�%I�D���}��Ψ��IS����x��₂TG��znV;Ll��73T�_�R�e�JOW���U��N���k�z��م5R��pݔ�c�=��>m}���n�t0���������}��q��� ��� ��I�@�k��k6�1�'bi�P���SC�x�$�ތ��L�@��$��3�ĉ�q=��Nx�tВ���m#rriPa�ıBS��à�����W1��%��u�t�mc�t��y_�|�#�C��t���a���!��g�!���ڕ���L��Z0�Z'��X�����EY���Ȋ��)_g��$�@P��=_:�45_���/�� �j�g�V�"~�����}D��Jj<xi�4�)ޱ~y�Uvnx�����wn�q��l-�9ʨ(�݃�,:3�8�MH3��'�RN�c�,�b}�wx�!�R�>�����֧�iŞT��?�?��A0`���K�^��L6�g��ۀ|ip����C�X�:5s��՘�Q	�0�8|�}���Z�C����:_K9L$S�C���IE�,d�V��6�j�&t���qWYZ��#J\�JK��Ph��~�svj*�tZUn@�B�.I(�2}ǲ�ڇ3|�5n'	�po���>qy��ɦ8ۖ�&���-H�?���
P�7�F;��8\�@>i?�k�.;�׷~��{�<r��,�W�0\S=XE�bB���,I	1��0T���"��꒒��8��_ ���4��z`�5ݨ6"h0o��Hh��Ƨ�2$�o �������K�5Ǟz)u�<�k#����r�ϖWbI�.f��E�j�0;���&�O�U��6�D'�n3{�h�*��6,k��p�{�M�P=�g-)\0iP���x����+D�"�1�Ukv�+��,�-������O�א-y/���=KWݓ[��C��O�v:D���ƔM6QvOˇt���&C}�T|#��9Fض�/ Lo���5����ͩ#He\�>�wm��^�
rб����~(5Z�1��K#���~;���Y�F�r� Ҙ�-�/��=t�1M*���=,�Vo��ُm5C͕5r�g�R�X:��0�@?Q *=�q�E��1����#]�����+}���*��J�k��>~�����w���7�ɚ� �~$0(��*EO��R��D�3/�+����������O��<��V�Co�Z�ZrJ5��Зp3�!���l��2e��dxy� �ޑ���`j@�A.C���Ӈ£ކcُW7�B���;�5�4��Uƾ��2��%ejb� ©�g&.�����ݘ���!`ϡ=����y�{�UWw_���{��� dn����tj�Cր֍-Zʛp�;�	�-m�2X���X�������j����lJ���\���a�?���I˸v��4�����^
@�]�jFߝn�q����!�3���R�%d1���3�-4%�,���s�	�z��'��o�/L�E��L5�p�=�����y�K[��L{����}t�\�9~�C)��%��-�k�5��Zw���K1�:���4�3^�(���<�0�D�_����H9�(y�!���%��H2R5gϐֹ�B�G�䀜���;>6" A�(�yV�G%�5s��ap/N���~IS�O�W��QBx�'�INB�z�U�Q�T�V\�(��o���:0�C�?�B��E�J�>ւ�[��o�b�Ezu��HE���,�w�;�K��Sk���2���ѝ<�Rp.�W]+=��s��e����@�X�E� �{��:w6c��A�q�qe����+~V� ڑ e�dZڪ��y�-�i}V:�L����h6��QW-`�@Jv��{Rf��N�,����A��������f���qD��ļH�Չ�y!tS�zب5b������K��E�@i+�of^�ZR.
�O��\��W�%JK^��f�۵��+����G{��H�-�X�B�X��$KV�G|G���̣$En_[��m@�z'�U2=���vT8�\���#T��c� ߳�j�9ˣru(d��/ѵ��n���Y�d�CP��Hr��9w�<
�*T�{rN���1�C�����7�tƦƲ������}���{���/�c3	���&�M@��t8��g����q�!(k[����'��{"���K���MWf���V��Ú6� �1�"���N�+��YKj�2�w�d��.������ՙ\�>�h6��`R�E���'��%h&іu��e�\vnSa�O�R�I���犑:�T*�M�m�g����W.a�3��)�S6�e��Q�KC|�lB�	{b����j柿qLο��+�1[�BcY����o�����g�$��&E��dme\����s��u��2�K�m�����m�g�x�CA��-����e��[��*d��xp�d�y�� ���'&�h���Q0搬x.'3�E?'O?9!M��Zɕ�kw\��M҈�W9Vēwkm�; ��������|��s���D���E�$It�[�gw�������5r�O3�i��ݹ1>�*P*��-�K���g+�� 2�����<����Ɣ©X��	�{�+K�l�4��#o;Dq�8�0�؎7a�y�ָ�g(X�Ș�ϧ�*��k��+�hP\c&6^D��~����`�4�$[��I(�ʛ�x�,�����cVĲP�Y�k��pI���e�P�6@'�}"V��Q��x�j�}K�P[���� �m�`�{�ʛ=�cu��i�0�]Ko�=�[���w������9%����+���l�Uca	���{�� ~+�,��^0�I��D�dz�W~C��D/��fz��$'9��-�{�i��ǝ�����GQ=�����sZ
Z9�\�7��%����II�v-���,.��V	~YlY΀��1�@7HԼ�c��w����x#��,mѪ	E�U�S��g���H)[�Ns���RK�_�}VY������T�՞r1W�֑����� �M�{j4�;X�¥@�^r�}�k���K����؎<o�,�zS����sr:,�!Զ���o��Z^ϥ!ױ�� 9X8l���š]��[u�a7*26Z. ��p�m{�s����7'��ө��d$�fZE/��Gm�T%�����0������^��"�[QMDmC.�g�G��+��tcRKJ���9k��ZB�e)3���:��b�D�֝�tM�Fֻ�M#Uu�LK�4���;hr7��z�On��I���X/
��Zf�Q����C�u�0g�NV�;�YHa��ñ׵>���jd�5l?���|$���{��W��5u���: �"Z#7�ҋ�+����>�X:������~�s�	��B�p辝�꧱2�ō'@�+�9���&�r���Ƽ8�����=�h@��k�9H�іz��H��8 �(��
�K�ʏ��@����Qxg����+-f�d�e_9%5k����O�g�N�A!�k��5ن�,L��t�(R�~��8��֝z��֜a�N4��ݥ*�WM�&�_'
f�#�h}>-�C@:vǦ�TPeo�&P 6�A��YS�jt�|d\p�y+(�O���3�r.����	H�iKf�F�����y�l�a��d
Rg��՗�L�%�T�E�8�B��*��z�U��3�'���<0Q�,��fB�-�~B�B3�#A]4c�Q��; ����s;V���2���F����]p�1��|:�m���fN'��΅vT6�3��BA'�yq�j�=9z�y����n�+/��}���h�q���}-�c��/}���>i��A�,�lP��N��t�W�y���0m���� m�� q0��S7AD��V6���>���^���ȡ����*�ݝw�߈����	�N�`�ݮ�
���mwR���d~i���d��z�o�������^H'�Q��;��e�x���� �Y7� _6
����+9-u��&�P#Sqk>���E�R�:��.�Ӥ�Kd�(�k�� �𺧍�V1w�e���ڒr4|5�V� Qo�����AIHѨ{N)D�E$���5p4r`�ۄ���l�6��fø�X��{oE���6���s2��\�S[�k2�~Ӧ��0�w��ŀ�j=+�SJ���B�-Icz;�߲�#`�ӱ�3l,X�H-��G�:����δ�Z){a,�C��Ğ�˜��?�e�o�����b��=����>|5<AY�	{��37�F�2!��I<К�5?�IT|����r�K��\ �	���RE�f�&��-:��5�Gzś�--|֥=j�v�g\_�����7�L�Ϟ��cz���H?��QL,W�:XӰ��ĤI��[�=0� 7b��hD�8�
����L����r�����KD���Z��&�t6ڞ�.���x*P@�}�tT����D���1��ҿn�_`
�޹�(�U�K�Fp���P�e���'m�G_�Z2�j������G���ǰԼq _c��X�����/��1&0U4ݲ��2(j��^�����)������$6����|�[9CƝ�z�^=a�K��tf��e�*wZj^��7+O@� �*[�OK��t�GE+N�X|�I��$��ʽц�C��є�ܴW�P�`,{�C5�����@�f�B�8�H"�==�P���/��A>�+�837霣�k�,
�63��P�Hy#�m�np�V����X�`c����Uv�᪪�#Lf�x�"��G�AD�r��R��}|��p<��S$��� }�;�]�ڜ�+k�_�E'\{p/tw���B��@
��c�=Y
Ȭ>�z4�LX�4���+*�O�'�������/a ��X���1٩_��0�����+��||�a!$�:Ω�J���,B?36+�w�C9/���	�T;0�>�] |Z��R�<�
���<������)�~���.�Gk���!����a8��_�����8V�b'ײ@pk*wh<��v��ҼU��&���)$������/�剣��ľ/ػ��!ZFv���f���b2E�}D*Y�����'mG:E�"���[���I�O�#x��u��> é�*C���M�4�%�c-H�N����4�TAZ1���Y���Q��zm�95V��>�2ߝ|6N�ǔT�Xʹ�˄6�2Af_g\��i�@�[���ˎ��S:�	"A��L"��(�����h�|c�%?�}��4�QeY�����aa%<����8*�P�C��rb]���Ѳ�$����Ux��LPG�`\�m����#��Ks����p�z��6���BBV`����934�����RM��6jIK�@<��q&MI'ٵ8cr�Wg,IXb�G� ah H�X
Q�=1�:�č��MB����Mm l����+������\3��#a�7��R�8�44�l��=����团Ã~�Q���؂0ܰh>K��s�ok�>�w���\ܽ�M!$�ӫ0b.����4~��|U���|�؇|��H�(^�����m�,�y�����yr�<hn4W�E�J��g�h�Ѭŏ �ͤ���'IDܣ�Wn�%�ݚe�(�*)8qYds��27zfB`D~��pb�5�8�ʥ�@�o���+z�;� ��-����oӬn��{9z|��g��C��3�&�op��.ܩ�iW�d�(��1���z�GC��<	w�	���5�U� �2�L��^#�&�T�r���a�Ⱥ��$��������?G�E+�V�V��	��~c�o9��{�꤫X����J�{��X�
�etV�m�+�:�Ԅ&>�|�AS)Lﺏ*})Ѿ����t�iR��rzc�~����6�Ծ��AGb��,�SE�V���4r]��������K8;� 0-d���D:G8��T���u^KX4�.��;��j�+P�R�޻-Q��1�R ��n�QorE�*����#�WX�����7~fu�Z�����H�L�E��LA��b��"��I����#RS ��O	|�����LDx�+!�6���VD���%!���GiM�t�<��:�1�ڭ�13�5����������'/3��~S��o.^�� Gļnr�W=7Z��H��BT��#E�]2�&��/��,�o�(eV.�<����S�ε�aл*��fߎ�>	��C��B��8*]7�|3$�Q��m��K�r	�j��Rn[������� ��L�-��DEq�����2~36.:V�����'4w�C 9�����O�C�q���Xx�z�p�QĖ������)c�˯�s��Q�2��j��(H���L��{i�M;�,��0ϝ鐐V*a����&5ߙr'����	�&��0���{h!^]�A���KK�l҆C���vA�+�����KB�F��<qS��f����̐.��G�2�z؁������M�K͑�ݣU#�ŻӃD�[q�y����BR�ԇ2D��,���ð�h̢�L���f�~	�W��H!���T�/:�WG��NGjœ��o����:�H�b8��SF`�O1F��J����O�S��r��ԋqT��`�z�U�ӆ�=�����\f?xq	�����
�ԱrxI�H�U6��S7��� C����O�-��Z�t1�m�/ݾ��5��mɠv5v�����O�Z��z�<���8U}��6e���Cv��庱*�V�`�k�K��xZ���+6|USf0_Z��цu̴���r��5��c��=h�$$����~�7�M��ΒR=e�Ѓ2_���q&x�=�΅�0nD2:�x2��ۓ8v�7dD�J��H���`��j7�MmkګZ-Ȁ�I�O-$��9�pv'�CeZ7Y�Yw;�	�Ul��Dfl�Me���AN�ִ�/����,�C$΍(fW�0�Iv�&��({�l�i,�Qru��A���\��P��ylD�l���wVn�KbA�/n�';9v�xǑ��D)1(�Ue�0��3ЏRc�{%���Ent������*����T���X�� ����KcڶY��Ų����s��p�K�VP�����İ2t����1�ǌJ���vw?X����q9Z���4LB�t��uV.���I�[�zHO=�d���x���F�`��>�DN����� Ű(��|�VAN֕��_�5�kcj�i�ʍ5C��&.��*�jG����_r=w�*��e@��U��gܝz�E�,�5�ܮ̟S��;���_U[M�#��S���e�[R�cA����~?+��"f{bC�:�����&�P�[�.�z/��Ƹ'2,^0�6����o�:|�;mC�(��lr�yж���fa�^�\�* ��w�U���Yd�?L����nBK{J�R�P�Y2fѭK�*��B5ġe�d����븋��IT5�j40,f�W7�0r�|Irw��rK�����A�n�U���>����DT��V��5D뷒���ws�Ŏ���~���Iߥ�pD�NF�=����Q,���-���a ��/�g�2��I���ap��zazm���0�w\w&p�����T�q��OϡE(´q�}�eKV#�5�H�=�N;���4��x�l�`ü�Q��Z�d�p5�.�_����8��S�x��r-i;��fSGt���p^�n�N���8U���<�2J��+Jkwz���fao��=�g���7��k?�_F_7���rb�лc}v}�?�����X�(G�OOS��"P��sz?�������9
6�r�R�0�/߳���7�l�H��ـ���D�6\��>G#�����@u��a9faP_�80��l�=�&\�d���'Vt�|�t}�+���v-��-�&^�@`z��d�Fa�����;���X�X�Y�Y��^NfN�W���)��QAE���i��������-k�O����*uj����#}}��O�p�h��;�˞�҂`Z>oHL��x~z��G2J��1���)�	�D|�2�k()��bM��v�muz�cW���b��S��*5i8�+,;��S3{s�U��E�ٲ��"#�"{�Ri�x��9IQw�(��VF�\_)؊w���+�}��t�7�L6�p34Kd�1�σUP�TW^��ؖL�=�򯯄������,'#%�r�U?��A���I%����x�_#'UNE0��IjD'CZ\���=!y*pdh�1�W+`2o���Z����é��`���f���s��A�[�8@�{ۥ��vI��+���B�f�l��.N���c1�RT4�v���Q���S�c�a2�CD�;��9��~���bM(�pM�@[S�\�>��U�Ť7'�l(��㙵�����aO��bۡ:�&�As��I����m�N�gٝ �_K����eZ�b	�z�r�'���ZB��uc�lHr�%���oj��L�7S��1�f�!�� ������z�r�ا�: � |�6��N� _��,�N.J�I���k^�t�1;/��&K����p�c��^�s>?p����4rҨ6Fp�T���~!����� )Vh�)�檕�"�<��tsqu�w<<PwAx�?I��{ɉ�8�c�Z�jXJ�=�mO�,��v�Tٟ�ӻ�[Oz�V�V�/�&��Hs�G�KaܡVo��#4~��,�-��﯎_	�|\*��k�<��=��̴����1\ı�x��MZ�4Q�xD|��vB�J[��}q�
2���k�0�Q�>/'���-�;M=����$�bLr뻫�������&��S�8M9�ϯ�4�T�]�땼d������zY��
 �l	p��0���F��rQ�� �uF���A�6��Pp�V�t`0F�ļ��� ���U֧��Q��{�7(<uRf�Ģ#�V����sA͍j�� ��	TJ_�"�&�չ�r1G����!�d8D�v=�$^�ll���� ��UHuV�u��Y�a�{�zE������m�{�q��dC��N�^C(y�X��V��C��W��jO�t��R0^E��C��8�0��۫����V�fY�q�@��%��k�f���?R����G��Ӏ��0`'��t�3[ug9[t��>��
��գ����Y�Pj*q0�P4���-b_ux+� La�l����=D*�Xr ��� G)P��HT2���!m�� F� �U�~��6�S~�D&0�+������2p*��fKM�0'�A��A(z��u��|��i�VPg����A�TћK����~�ǵl����[����2Ɂ�4NӔ����mqr���9O���9m��ƪ�`����2!�4��LMi ��2�C',8�u4fi�f�ۈ,gݝ:M�����Z[Qa%O��������i5�fi��/�|4�<�NY*�m�Z�t�#��'׌����߼�UA�.��zv�)���KQ㼌�E�!a	M��T���)�+J"7��η�>���~-�0��߰X���+a��������6��3K�4�6�2����&�#b녃���|��ֆ"?$��!�S�Kx�)��������{����2�n����i����E?�Z^_����&���p�f���O��^�C)�0�~�����O����2,��IAU,�3@�F�<��4mQ�uB��|ԖCn��c!�=�k�ݣ�� K��VԚ��q�1�y���p�#���!��Ϯ��	u��L*H�t�ꖇ
�k�$���p詥'�uyn��p習���H�EF���Z���I��=��L!H��W���f�!z������E"^��v�.�G�ڪ��Uבּ�M!��|5,"���Pt�$��������S��
�Hq���_/�f��#_I?_���i��[|;?���v"u�~3%�!��jI(�'IT0&�%���kU��y���B,����Q�s�;�[K�6*�!��GjD+4<�]i�
�ذ�@+������tg��p�<�c)��6SO+������Oi?�����+�9"�vߨ'Wj�iۉZ{���~�LjH��Օ���,uV�T��T�e���K\gy��x��cy`��s��d'z�	�ԋ��@U�<X�=��̃p)�X����Q�M#w�����E���ۢ�P��ʊru<�(jd��C�7"�x�@���G��|Zr�������vj1��`Z�@�K�������1#p}�M�������0��k�׍]0�M�J�&*�[���f�4�[U�0"y0�.�+�k�D��դ��6�o_Ez�� ���_��L)�8��8@a�T!yP��N4�O��I���;P(��J���:�u>y+�N��w��d�
.���}LԬm@2U�³.ITQRX�z�}�\�W��)�'�g(8���kN#`�Ri6��Q��H7�a��<Z��=^]�tߤ�Wnu�ԅ���V5�U�E��P�(EЙg	�s>��ٌP&іB�Q(lz�z��.��������a�/����yoy9&�� ����v�o���٧��>e�{�h��C��t�� r��~.�,|XO�s�%���q��L��䋈92���A�j�w1�Zq�,99��Cy0E�R���D��ݴ���b����W~R%ݿ O���K��ҿB��t佔�q��Y�[D��k�6����v�\���v���ǘ���(���E)�ܱR�n��1D���sn����2�SZ	J��?�;�N#���.4ж���Ȝ�i=�в)��!ᄗ�>pA���7h��(��ןe���GG�8m|�����Mot���+Q�:�I���g6+^�g3c��?G�w!���j�n/���u�
���d��ZvH"�>�������%촉7a�P�P��J�j!��}Aѫ��3=r���<pY�YG �������%keL����?������<��$�Ԙ�*d@@�=�JD��+Rn��Jy��R��iG�O���|��z$eP�# I�DߑE&`\�K���c>�K�~��UQ��%B_٨)S�B��) �uB]֒8")#b���E��R�fƼ�)�ʥ��g��-�ksj��s�PN/��L��]1��3�O K!q-E/������x2L&p��I
�]�Z��5QK#�Z��DԻ�l�E@���v��S�v����� �#��}Gτ'��Y�nV�%�᢮bh�wT~$�_��AF��儼%Ж�*����}��mT?:��I"�,���"�޼O�S��?�ߢs�IH���4~L�Yh΂w��Z�X��Z�d�չ�!g=gc�d`��ʃ&�tdlՑ�{�& ��| x��� �a� �ֽh��qE����j�5�~4s����� �U�r��E���Ͻ��!;�9_�.I�Hw/�=�D�%�F������tB��v1�@��� 3�ֱ�E^��	��?��h��"[��s�$۹�B������u�ѓ���^\�)�}s��Qa_[Ji���,w�<شZ_��p�ר�F�;��)z��i�Xj<V�"�尒������� ��>0H6�$P1{�C�D$b47}��4�~��AֵB�Ҫ�vGV>���kՐc"?�X���@�6��Y-�G4�p�-��zp�Q?].,�����Q��ޜ���(��L�Xz���M/��iX��vD�N�P�
�l>5�O�kå� �+)�|y((
�O�,���o)^8�mJ�ݘ���t�8�S@Q��jݓ�o��ƪ��F0��<�oM�4�=g�p�����9��I[���Hɖ)w��ӨF?e�;��7e8���N�|���̀˹J���F������x.��n�@6����0�D��Ĕ�Ƥ�j�Hr}�P(,�#��܎��V�DJJZ�Ҏ�w�*�>tU�_�A��V�nO$��N��L\2�4D�`"�'�$����Ι�[�yI�Mvc�	�-����w߂�gwF[�ag���`.��0ʡC5K�Q4C���]�@3���菭�H1c��${>	���]��a����_����Iq��ƫS���"�&#��≽T8�3&&q;�� ��-�=҉��9%1`�n�G���� ��Ϭ�Te��&Und.�*ί�t�����mg�ŗ��$���A�B�o�h�<1\�XF�����7-��I�$)`���Z1V����T]�(0Լ��v�6?��z�c��/�1�����wb4�tI{_$yE��a�u�r5`)ڀ��7���	�4.lX3d�� J#��G��栫�1�ed]SU�ħ>��(��6���l�\��xo����Q��<��$�9k'���{��q���U���W���z��=��	}5H=" �X덩������j�gJ|a(��M�TD(�I��en?JMZ�mH�g���i��b�(]�Y9�o�\	��d?��*��D�Q�7 �nGk�t�[H���F}P]SN��Isԩ�S/�W��]Ce5�D�J*st"RDqz��a�i9�fh�&�a
���)�k�� �~��#��#S�Z��il䈹X�lp<�t�����T��}��J��#9��A�Á���e![�e��	V�������P^ͱ2+M�s����	m�j��w�XC��TPS����P>a�a�ig�+��aB`�YSQ?^qO�}���4kE�_|�|�t�|���05v����M�ǉ1e �c1h�+����mܞp�j0@�	#���j��.N�I��M�hc�#���|��=���_�)�k�u�랅��K�1T���˹���faZBa�����Z��ۙ�ި�5���3A.)�^�>�#1�5r��)����{κ��	����=6j���s�A�������YAS��a̴pX����QZy�#����� �X�`G*&8g�/@��d�}����xF���n]w� �����ڃ�GQS��q��^v@���t�}��눋���ڔ���?Z\��^$�}`d�>Fĕs:� bB:����l(�Mq۷�Ԭ��p#��T�D�<����͍��4��h�͔��FC��(#�c	�O��*W�WZ#�e@��qc�n�,)�%��~��xgh�4�����>�w+����[)7z�,��?�f���l�R$p(.���H]��B>�^�P�y��é
���IC, ,V#gb�\�m(����Sz�!��b �^��TӬ�O�*��@�8���@�5��a'�S�`��/�3���J�onL���G|RM�޵&��0n	t}�Bf�kh�\r+	}�{.�Y2��ɓиȾ��v� %Z�&j	Dهn��Ց=�H���<R�d�m�������@"!|�.�,oM��Q��Tp�b}����iYEe��^ޣkO�Eq�?����,�x�tb����@�P�ϴ���	{NQ{H�L#D-W7����u��|�/+M���Ͷ\��`����y�����Z{~�.�
>�׵&�t�MFM_/L_Y=��Zy�K��7r�
�lmBc�P'Y^z=��>���C���&�@���ހ�}lv<��_�����^���Wk� 4��O���D׈�=��3)��H}�?r��Y�J��	{�� ��O� �`��L�>��*�{ɔ͑��=��O���"T��&��٤�g�\�F���m��V!�M�"������X�+($�d@��q�U�B@�NB�3^��G8	N�� �!��+��^#�+[l�n�B�Bg�y�o�U�W����3�eS\?�>/,��DbO�9��E��y�g�ܹ�j@(��:�Q�J�w���c�ͣ��)Zz�ᄝ�gƍ��ü �2�1�_LTW!�2�R׸�I}A@��^�|lU�!.���?�ᶂ�R�7,�r�Ud(��Y^e�Op_��8�8��|�A|��H�yO�����y�2Nd��ԑ��B�t&΃��`S}���&n���O�*��*<�u���P����ǓKB�xt��C�3����Jg�՞��Y������A)ބ���s��2e�Uw����v�J�����P(��{EĘ�d#uDG�WIN�eIN�-?�Hr�j��-���K3�0���������b1u�yVn�?n�.=�4f�)�DMJv�W��G�����QV����.XE�ZUP�$`���	>���Me�9�U>�	i/��D�=�{e�w�y-���7j�
/�80�ʨ43��*��o���N�lr����誟hP��ԓXkU�t��f8E� T�&��>�e1�+����	�(���5�e��@*�Z��d�+駃�r���5�G�?5�'��o��j�M�n"?������n�;��8���.9��0��9��	�P�P+��Ԗ��]O�+�N`eS�"݋=F����S�` \yG�m�q�H���pvC�ᢅ�N ��p˱j��M�K.�V� H�%��[֣�o(�;F��g�;���22U���������3���*�tO�㤱���9%x!ܺS�����b{�w_�A��t(�d�D�ņ #1�LaR��җ1����M�t6򊛝�����uV�VĺIvtYSe�,�n6Gq�c�uA)O�ަf�9 ��[�&�i�[��T�~__��,���G����ű��S��o�1����阎(���!4�.v�1˳��� �?[�eY�Dc0�뱆��]�ϝv�;^]�0����][5j���L o؃�J����e�����N�o@.�N�ɠ�WՖ&֕G��MuT�QL;�JX�a|;ق,�B5�F��H�j���P��Hf},��Ob�qm�>[� gy�a��n�(3Ϥ��<ýL�Jj�ɏM'DͤeN������A���"	��l�ԕ3�)��%x`<��C��d�M��(�~2���$��I�mk0^����a�ؐ�ǹ;\-V�y��q��Ȗ�fΉ����XP}
:6�v�JK�E��0v���	os�=�3}�Gٖ�Η8�ޣ�7�ES,�~��$�[ңjᔉ�trmT���~�=�;�y��Ցr�J���z��}��鐵���K=������:�we����N��Od��Ìp����V�{�,A�
��Z��tL-�0M���Pާ�b�
\;�i��T��U,ùC�X����UA���n#�^��e �[��xG��4a�/��z���O
G�Y�fx�=h�� � m���s��(Ȥ ]�9�@��<��{Q���b�>@��Z�M�65v2c�_1���]DT��OkE���~u�U�g���z��vAE���W.��@��d9I�Kj�EdLq<� ̓^ꡮ˟&K`�����w���BZ�!"�փZV���{~�����)�u�׼��@�qG�x�QwxMr������X�s/Fd���	�o�\�?��(%e@x���L���g�c�&��ʑd�A/��pr��%����
�Y���T����40��� ~�{;p�P����[�;v���0�0͔�]*�U�F�"t#�f����'�V���"2���k���4G����$�m>���k0k#V�Ԫ��?܍�*����oq�v�ՇU����sޑQT%'�f�.?��\}���q�QfW2J���w)�c������c��{��g��^��eY�Ʀ&�-�� Z^հ+&�v8�BL�.X����\��y�ޝ~3(�t��F������ѽ�8�����#XH��.M�W��"�6 X�o���E�b��״y�������/��׏X�u�?N�$W�f|��|O���	Q=�M����/�n��A�q;/\�|C��� _�~�Pˌ�տ�TΑ�E+�]�~i�o�$�.�Ɗ��4/)p�tOZ�� O-@
Y؋��(���Z�IJ�C�ː�k���t�,�S|U�������v��n� F�L�U�5������m��0P�ґ^1�D��mW�0	�3��ꈰ��"C:L�˵�ta>�Fe�+�!U�F��2���y�$��Dx�5���X�<����E�r��%�:>�j�yn���(v+�"�1�\���;wښ��{�f�It5=�-)��dV��1�J����W5��YK�%�X�M�p*�
�a��(@�����ke�nz�]�*̢kM���/8uǳZX�
G��c@
��Y��X;�6_��q� �V����+�~O.�Z]
��n�~v6?p�{3��ٟ�H6�#2�!Gx_UI��%��&X���+`E��@���xaW,�b>����iv�О:���Խ��$O;x'�x���Ԇ���^��I����0��?��4�0|� 6?:j�
��>οo�@!�j9�-LG�����>��6 ���3 ��20�7���������y�TOk�p�V������W��>�O������@�	�x�.`+
~�������y�ۭ��+Y�ʘ��2Ҫf俈^�A|��^Sb���%�,-��-=��O�'w�\]S�.���P?o�`� �
�~I
�����G��`����M�@]P��w�*|��4�["���2\O/��ɶ�?�=θ�~[87�6��Y�V�h�!p]j�;���5��/�m��1g�a�l��4T ��R1�V3MEB�,3@�$���kh�`Ϣ^WPl�����	�rԑq�Mah?��i�
ڍ����Gq�$߀BY�{�}�兕W��`����y_�l1�^A�o��-1���Bs�w���ԓ?z UU����4����V���Ht*'�Ž(}7.�-n�q�#�ɞ7��yv1�����w���C�
��J�)t��w�v�T@n�.�VBt��;wI���Z�����4rr���0��X��t���3�^!��9�֤�f��i-�b%�ޮ2v�� oV���Z9tC�z��s/݇�#oÛ萬�����q)+!��{MBO��T� Mè�:XI�͍-�������Ҋ��p ��P�t�9�駠եpl��:�,R��+��n�N��'�>Z̫eU�,U�����界��ɿ�m)-���\{T|����ނN�}�PDIbT�6���RvE�����]���|�0�ٜ(@al������x;)fn�⿯���ɟU=sOn��B�Ro�lc��E�Ib*��e���6,���yf����k{�{�j��F�����Эw�!�ӿ7S�z��q��QP�Q^P2���I� �H�߫h���=�"	=��ƃ�D2�W.�Xo��Է�&����
��9h�!�c�@�w����D�'gTX��?���ɯD`4�����x�"���MY��}s�d�Ɇ��ӓ��������2�\\��F��,���k$r,��+���A]�,�((���U(N�%��ע�
7� �P��"o�^��Jb�^�8���Q���eџ�z��@7�3�*��jM���+�:$��-�Q;D��@����QN����v��UCm-�v�*���,g�ҚA�M[��F�����)0e&~��A�dX'�����^��a����u���5¸?/��GSc���씕?K	'x�Jr���m�ͩh�E��-�i�"���� y�U��?�
�1w&����bQ����B���y���,>��s&�)YGj�bv�r&��P�RâC�dhsde'�5�tGv,��sX6E��т��Z���3�&�y�h���#�%B�I+1��I�f|(j�Z��LՂq�K�@m�xxŲ6�"����b^b?�������N�H�I2���?�p�x"Z�z`u�N�����d���(����Α1qi��K��׶ N�u5} �W?p�C��{��."S�s���H��O|6�~�L�d�/Z@u��#��0�؋���\����$'X����ak� $Z(�	���Cn��o$��d����2�eo�� Q���
�<J�xh#��cb<���{�.�����hɈ��Auܚ����|X�$X�<���W�+;�.�C�X�{��
M��C<���4ΒB����~�|��	�W_�I�3�*�lj���3e+ٟ���]%LR%r�@I��R)�*�[�%h��O�I�`D�7����gn��aQ�!�[��z�I��-�域�?��8-�~�"��Y�E��(�J�"`O��Xáe�
O���s��p�f�J�������B�B�����K��/���-�e���J'�-����!�D�Gh<���n��z�Ui�d�����D�����|�8)�K
��=��
.
;g���7$�B�	�+��:�A�Ki�!D�9�E?���ۤ+�ף�V�$&�v�@w��^G���-c���#��^�w������/�M�Lisl�{�UǠ��+�]�Ī�딖e� �=V_�Z�o�R����y��rG�ɗ��I]�G���cҷnQ,��~��]�npi���%��L��-��5I"�7B����>U�c��;@�`�v�X�X}���K��ʮKq3� �j��I�F'tG�,��[?��z�������=��k�
^`v��E��jG0t�|F�_=�T'-zeØ�����������K�;�G��/&K����LQ��:fio2��!� ���7����}��~�5}��QCF��U�?�9D+���cdcn[#�s��6��B	LRDsj�����;B��Tp�b��Y�<��9x�+��"�x�����):!�+g׎K͎t\���^��	W��ڰ�R��y|���~�㦧!G��K������#Ǟ�]��l-����W�"�)��6�ौ@?�ɻ��a5����[b���i����V`�� 	H�!�^�$<�o����J�V�2��r<dc�6"p0�2PGG"�J��
F��9�ᅵ�Z��
�Q!�8�w5	�q��-*����ɐiS��B[�1�]5oD�m��`gL_��?��+�ܩj���l���]a���M���Y߀h�XQ}F��v��㮫��8�C�v-C��_���I{}�(|�1�l�E�aSլ̃��EXT�N-����!=`v'�k�Ƒ���E�x�8�_�XZ�#V�F�üm롟l������ڊ+1�Wi��߰	�L���`Z/�F�mWS����(��soY�v���a�^������)�LVo���E`�!�tg�����P��EM�3�M����?dԒ���z�]֭@z1�৙�!��`�[+tN��2��}@��(��,�����H�+���?LQ�ݠF����੔��5׉�*#���N�t4����KN,0����@1Y��d�ܕ�=��x��e��? ���ǡ9f�C�3O�R���`���7�B1��~��ir/��������b 2M��<h�R����˔7��i�	���2*�G�&pW����j�K ��C�/��!��L+Akz�wۙ�Lɡ 2`ց�Y5M�2���4\�ј��O�$:U�ܑ����ٟ	�[L��ʎ�z �g�����Є{;Jnj>�Ϣ�����O�#l\yK,�sC��W-�%��U�7�4�yc�Q뜏�T��W�6=���c,j��F���uoeWZB����*|���*.����'���	��	pY�DS����ġ��!X�s�?�= H�twB`^�V���pA���W�:��q�m���l�*	^��b�P�Rs�@���}\L`�$���h�i�	q#
 ��j�/j�i��<M��YA3M.��K��$HL�^#���,�~� �(���*z�]��GeD��4P
�Dj��+a���v��Yt���(|��������ܞ��g�A���k��b�W��ٝp�#�w?��=�/�K�OT��u/Nz�%6p=�O1N��^>(z���CNez�:���7�h�t�JDG���d�BR�����^�ª�)y���"3Qlh0v�t��x\m�;�Xز7�a''�i��c.*[�]�E��b(Zܰ��_��9x>�'��
Cٖ�,&�6؏��>�~�0��v.�� 2��] M��tT��kĄGv1E���4+\}/�i2dK�?��.�]�/,�Wo�bI����jȡB�#�\��E���o��`������8JI���
����&�\GP��ל��?��s��q����!�`BqV����> �|��^��5d�`f���d�oX���Z�CLf�y��=	S��:����-_Z��x0�F�hL�N-�=lX^���9n�'&�5F���^����	6��Xy����=��X%��55��
�|�?=om�� ���A��wN%��Q��l�W��a�x)'�	�h������w�"�م�?��0&�*��!���z���!=��jT3z:�����#{������)�DEp�yL�-\����GDII�z�&%sX�����0�M��L8T�0���i;�9q�E<k�pvUǲ�˵%��m��X?s�YwK��ֶ���2��Dt|��~�r�����͑���>�6�4����R�.�������A	�0�����e��Idɴ�h'J昝�'�'����W�������$�9��|�UF�~�X�Vɒ��/'�p��|���ft.����mu�Ps]����վ�B��b�<��۱7\.z���j�L_�P!��N�fg���Cu� ��-d��DupҠ���T��nRtޜVb?���ˋQ����tJ�O�'X�d�:�Qq��pz���0�vUW$��֦H����l`_��Qr��y��V��J�Ds�y��t�޲��:��f�j4���P�B���J��]�-:vR��cpot��f�[��e ���FlJd|�9�����kj0L�f�GS[;���%Һ����(�^�ZJ�1!u�����&���[�I,5U����>]aO�9U�t�K���w�谸käRe� ��6�M���2��:B�9ë�nJ��=�Y�P�Y-��{B����>0��G?u,ݓ�e�_��í�����e���D(�;? 5�2�	E�n�Z���F�ﶱ)Su����5��_�L�,�L����T���l� �uB��q>B���ޢ3�L�=9/sqa��\	Yli� :W���
���*k�C.I��3��El3K�l%��<��T�lf�膫���*�Z��u���P�c�Tz���E�&l������;A�%E��W�f��8	@�r�B����͇=<��`-�����"U7�^�)��^I`��,#ܲ�y��CW]z�7UO1`i<����_�n� ��kwZH}�0y[���N��ra��	S��<��#�V�uBP2P��s�Gɥ�<7~��jm�$�8[��Ip��j6]E�G�^�h�`�c����!*3�2�>�-z,vEMҷ��Hr��BYh��<:��=�D<�>׺�j�{���'�,N�]�Ͼ�VfDQw�H���m�2�]Hh%�
�39�@�&)��CV��]��.'������~�-6�N�іK;5��ָ�I�D��N�B�����'� |v����n���Ыtz!ߐ%��冱ƍ�Z�|!��b}b=��M��mȕݒ}O$@ҔO�=J?��H�cď���?T7s,���aS���Z[CvTʋEA}�-�����h�HL����>o����`yװ�rT��(�6��w1�����&o��J�UՂi�#m|�5*�өW�/��d�J=ns=�
�D�;�)`u�?~6~
�M�]�NGg��s�
V~�hI�&+��=#"���� Y��=:Tt���^现���Ϩ�*v<���Y�y}U~\���!��t;���2��ӥ�0I����7g�a�=ٻ��Y��B��e��������^�y<+6tW���&����<�}XT��d���1$A� DjpZ�°���=���K��$PC�}�٨�9��)
7)����`5�J�2S-���U��q���J]#o_?�*���J(��8�s�mA�5����}��/�X���q�/��d�x�Uʸ�?��K���pl��$���W}�I��Y�֟�������k"�I;���|�s��I-Q�{'�YڕУ���6��=x���}-0	�x#�o��͔��U�P��,�(�HuW��De�3�p|��	1�J�P�E/S��(�Z��_� o��'J��z��f�9�]ha���q�Z;>�R��苠ވ��P&��>���Ӈ����R���Z�0��4T�����3O����Dwʪʡ�2���pJގ�INYA����+��_��[U�o��m��ЄbF�x�� '��Ҍ!8�����-�h8�?�]���F)i�9OӬ+څ�Y���3��j;%���dz��ف����k���y)%��(Rb�Z�`[ǩx�;fA�,��/8P(A|қy���j�Z� @��Y�}�?��ui�P����u�?k����B��MH)��؍�'���rv��$s�����y��*�d�����7V�m��<��@���wA.�o�R���*����.^��!�d���0D��dD��lY��ǩ-���5�n�[`�ǺBA&�eP��U��6s|�n�@[�^f�dG�"�SȮ_�CG+�������9;D�;���W��ժ�.��1m����&e���
۳Z�Dm Ad��S&�Ui�b&ߠ�Ʉ�a�	^�鼤��&)Oө~lT����V=�p�#%����&���?�H���h�!w;UC��
����j�M��ʷ�`�<m�\�pr�}�W�ʽ��敮����̆'�� am�-��~S�N)�$H?~Q��B��N �	�>\²�,�A����@�0R�L�B}tr!���吐��B5��X׌}�!����D������vnb��¤�D/U=*�I��B��ȧ�c���|2fh�Y��8��V�:0��ny/��w[o������!P<1;�m-$�A}�����!��t3�S��k��Ȇ�&�6~�PƖB��2e�:��^<)Oj�
�؍k+y��>m]MJ��a
lҦ|��abN��ѐsO+�DuK ^�/�!T�ie��%|�f�O���M|��n���'����+�$ڈ�?��WgH��q�8.�_5��� �,>if�g�0}�����Q�^���]D�d�6_��;G�6E��M�ǉ�%}9F_���T�fr��Z�Wg
���r���(M���P,*'��Y��A���湝�N�.ߨ�|;?ĩ�f J|kaX�p���Q�j�0��Yl���{��� 	��=��3�k�F�	�JE.4N=wFJ��:e�B;ߕ`�k�M��V$n���~�;ᔜ�]3���2{��j�W�Eb�Y<m*��"������`����/?
�%Ġ��R��I����t��luP�< ^NfȺA+i�cc��"V~I���ެqA������_x&{�&G�[)^��=�I%5�{La���.�3"������pb�տ#�$gU�<��ؼ5L紮�L�~�n�n�>�s�4
�ݻ�P����d�R�u��O9CǘF�ir��`��Q�6:�ƹj�7Q� ���
:�Py$������T$t�C�b�����(e���V�a`���(?k���#agk�  ����S,]�Ԕ�{FJ-�O�ߩ��,�"R�NGY툒�L>��Z���i�M��<s�}].�r��ٜ#2�Pb��r�c3������W�x(j
B���+���Q�׻S3�n�r�<z���6W}�ʅb��y2��Gk��_{eY�B��*��?Ë�Rc�
q�g��%��g�Hb �3-�z]
��[r�H����ߍ	��,/���(����p�n91;熁���z�'�*,��~��"�g�}�.>u-/�GF�_���,��㪤�-Zے�~�-�< �sr$��9ʸ��(�n
u+fJ�i�>4v�xi�۝H}mj9:���%��j|��tx��4l�NKt�������t�`�t�Y�M�@y#?�_��2�e��ҵ��o���3�-�����Q�N�"�Cƚ�5�&~t��A�G���G�S�ې���,��~Wi���#$E--��N��HR�]�z\��B?��u���{iJ�ܔi�4�k�w�����V0�'�Ź����]gkv���;�$�t:�p\Ugv�<5z����\W>Pn�Y��  R�ABj�+� ����2J���1���F �J�z$F D��l2X�~��:�i��2H����W�#1^Yq=���c���m�c��ll�&�������צ���N|�6p@2Kҏ	t�b������J2`nԚ� �˽���zcaM�o�p>*w��>���P�c��6�0B�/X�� 2�2�>R3_u�1]I1:�!��_�t�F���X$S|]O=y	f�bg|���$����W�r\L��@���}�D�-]���vHf:�:P�Q>��C�B��S#qq��OO](d�����)���81��0=��:[�z�"#�1	D�UvW��TŴ,���X�o7�W:5��ㄲrx\�d1� ��b;	{T��h�.���r�KP^.*�6�%f��8�Y�X�y

_.�EE�2$�Z[�,'v%��L�*�Uv��H�Ht5PP�D��7��g������&F� w������F\ �qf��g�� �
!A9���jeKmt	��p�SC�7��^H�=�׭K`�4窗��
�O�����sl���,�O�Gg�ş�9,u��y�g���I�"ڣ��Ob�������uג���q�g���ϰFh��憭��J��i)�O�D��������2����
\C������R�U�ք8��K����+U�A#|���0+~�	K��:��o��(��`�"�:63}S��z�p~�2a5=����𯉮^[C�b����3p9	�S6�E
�k7�/N"6��G3��=g|m�����L|ϔI�8��j��(��M�G���+����������8�w���~We�n��D�&E^���#�A�����C�;(���Y����5o_�ڡ_�ل��Ϊ�L�lE��[��թ#b�@D̬��}�@t:���tH��y�oD`�.ekW���ޗ��7�8D�~���QDi��C�a
�d9�m��X<�����󏉾V��)��R����xqP)�#FrmY"��?��}�&T�4t2��}�)p��.|ӂ|����!��u�ux#�J����?-��3�7}G���JT��}��:J[�#?ʓ�9�|:���8�E|xX+,j�[,�\S�θ[�����'�B�0��y����:�F���f�|�H��ٕ#���;��fn[!1H��*��j	 ������6���Vp �>��}K���OX��Z�����Y<	>7�$��@{��zk\N�z7�J'd+����U��b�\?f҅��������z�`eY
^,2S�,EZ��yO&݈����D��k>�-±� �o%�ϓ�]�f.�7{��}���^Cn�a����1�>H��Vo��=-�!ٴ\wG�Z-D	?K����p������q�z_0��;�:���C���3��T�\���3��+/�4�$�!��@�{v-�`IT���	A'�P��n��gf����c 1��b��W�k6�\���sq#�8���F��ky�y�)�Vd�t}��"x
΍�2���ʿ�m*:��]� @�<����ô�R�z����2㘆�lrM$z3�<�1P	���"S4�E�@���~�kK���EB8���?#+E_q퀔[���������:�{>�6Ѻq:5ɓ�=����^����p�&n��Z%U���i(�~n�'V@m^[G�r�
�Bkk=�M�^���q6�?��M��iB:�K'�*���8e=�+��c���V�[IX���Hu��rb�pP����:��"�]m$��%q�H�~����n���7��������Q�t��g�Xno���U��Ϟ(L���^���:b貸�e���k��6=��~�o�ѩYxѷ=�	�:��8��/�3��,���*��N�Bo�AW�_�)bΈ&������)Y��n(����-c�Fk��!(\��l��ͤ��3Vf#!�sn�c 0o�SE\:����GU\�ALL���,A���dQT�`7�9���ua�f��	��&7�Y������V����c�cG��W�d�h|�ʰ���'�i	 r'�W�<���` M�����}��� ���ws):� 8�J�͡�B����#è_R�%B'�Ѡ������)Q�,�ȑ�S9���~wD�ዝ�_����7���T������&�5+���rf��sr�𦿳h���'eyǉ$I�.>��N�%ʶT�q�G0'��z�k�"�C�����ъΞ��j:�؆PS��������aw�y���>���v۴b����u(NH_�V��^ɺ��Ͼy���"�gfnM��<���tP_��X�sqҿ��B�vw�7�9�s�~UÍ+q88��؊��ir�P$���B�xh�GM��G݋ʂ+']��iD枕Z�:�� ��!}z��?ǥ����&�A��f�CI&��S��04����E��i��@���As�L�.��X`c.(3b*�����H��t����<0찕g�v��6��=����,5~z>Q3��j�K�`VӍ����.*�;=@���_m��ѐє�`��Mv�}ۍ�.w�Ep��\�Y�23�"ϑ�|��e���pͿ�{�r��T?�X���v�X�����('d��H���Z'��K�
��J���V�>G����?�q8	"g����zv�*�{Oڧ6h�X��`��V�B�~ �[PIs-넨��ç��'-���>}�QV	���n�ڑ��r��C+�LZ&J�ۖ���^�8�}]�;�N��z_3�D	���5)��D��,�O]�����>�]����1N((�o��WI"֍����Z���au��V� ����dR�C��eld���؍��
�<*��`��#�q��5�KL"{'/�/p-�7�7��3�4��ȉ��ռm����D��������Q��<9f7~�%� ze�\`�p7��K��,у"/���+UMT�R,h����4`�o�p��'�v��e;���8�.t�l���5Їa��.��6R��矾��qe���;��*��w�5�*�;��:Q�� ����c��g�H��ѣ3�4�E�鍔�x��N��g�t�g�
e�����״��l���x�j&��'��dM6K	��<v�����pM4�G�C�{hKr����K��/�7�sr]'��8�V�ӆ�l�s������M���4���\��R�.������,+�"������5���:�m���Ix4�������% P|�$�!9ԙ�ۦ�ߝ}?��mk�����s<')�o�om��������.�§����D��<����������k�L��)��ң{�r�? �w�р;�fJ���f%�߫-tAf{�mӀW�gYY���r觸T��Bwlmd�_Y�>d�S�t�����N�88�+m(1�ѵ���̫S �k��� O����މ)��ȑ�7b����J��]2�����&��M�	���Ղ�3�H�M���>v��MA�(���u ?�|2����C50P[�����ԓ�s%�lKh}�[��Vhzp�������f�.ܕw)�'"K2n�6����p�'x*��F0��
� �E��x�{)���.��-���r>%sG�t� "&�����1���mԬ�K���o��/dS'�ـ�������I�~,݇�cr���e��߈.��n�E{�,���|~�r���u:LR>|O�@�A�����h�l/B*��ۨp����pH�M��T�!�8�~�E��4�x��w���D���HG�]���o:�����^�� ���n�c[G?����!�p@=�_A�0T&�\N�yX���x"�����Գ����8�j��w��3�ks�e��X ������nۉ�e<Z���8N>.RYɅd����4�t�BI�-dU���@jy�����}�`��ɄX�O�.z���E��qR� ��S���5#8�:��M�����-�L��� �P}�N+��2���_��f�n���҆��D��50���;x�d�2��ֱ�#��M�$�eȶH{�/�|����Zy89���~}���T��~Hd�k���������C)��V(PuK�V�>
m.���I�+  �eC!�"���TA�2f�V%�(Wt��*�&ked�ӋwѸdgm��7�0�-��[���b0�Rb/}e�U�Vm��0o�t�K�Qĭ ��<P|ӡ�������/�%(L��5��hb7A��#T�R.��Ѱ��Ȕ���)�6�GI9c��ܼ�I�����4��
�\|���X�]J�5�����S�pi+�nM-H2��L�=,���	��,�э=�+�L�t6ʒ[#ԡ������7�q��i%ATBcY����Qu��������?�R�%"9��ȡrC��ۖ���
ju!�j��j����t�a�M��iOF��f�h�d��{b�
!��l=�A�Z"&-���u��dmLm���B8���^�� �B�=e�E�;�iNR��������+��u��fn�dz�T�.g�ߧ���8�,�w *�y�������k�l�d�������5*���U%�ѵ����	١t�ҡA�?�]���Z�5< �.�l��w�s���7.�2N˞�z�J|�2N�=� �XXT�o>��.-�빷��*Z��M�͑d��M���S�x4B�י��I�%@h�h��gly�"�BU�e��!bBUfY�
o�ݓ4�r�*��L��Sq�lq�.B��A���Q���q9ަ��o]�Ni�CIp��jكGO��*Kd��Lp�]�w����4z[p-�ɲ�h|Gth�������%��O�p��� N6�ɻ)W�uH�{��t�E[��U�/^X�����Ԩ��xR(�bad�T��SJU�N�v���I;��7��V��-w�����`|��"C��M��:�8�\��5��D�P�I�L�1�!���#B��U�o�eXF�.�y�/��6�vf���"�g���&w��l ��������{9�2&yd]����F�2:֫t�X���)���棇*Az��8�%���Ѡ}��%։�}���$�p�8�ZLS}&��h�S�hcJ_Zs�?[3�y�ₚdgT)�(�y�7h+(�1��V�f��ϛ�e��j%��\4ur����>��b'w��b�kMm�̛o�M9@��B����i�{m������&B����'/�z�����"��`���K���e��-oK�'E��
s�����E9G�́��Tay�+dw3+ٵ,l��AC�Oʂ�a"�~}x���֚������ω�y�Lb�3]��7J���Y�]�@�����ZG��o�)(<G�FqJ��H<�i	-�dR/]��^��]��=����gD��ޣ���B"�Cş|��=H�;���] �J*��qx���y�I�Q�mB�Y9��Y��0ܑ�"��R�Z��@�#h-#�_VH�s�VF_�LV�Aׯ���z�g�V̿�_K�[�+j����dU+�x0�o/Yb����T�$n)~B����
�s<��@P��5=k�<C��x3;VS)h/q-gמ����n��F��J,��^zH��P�\�.Qn�:�mK
j��?��*M�����=��.G�*#HD����M!5a�����n��ٿ?��Ӎ�N��E�a��g���cw�!�Δ��,��s�w��TrD�z��L�����Z��)E\�"�X��6��=6�_�;Y�E����J�7�l*�������H��cg�q!���H���S͘׊~�
��ܳTgӇ�����ķb���SqIĶ����N[F��%3�h��Ι�m)2�������<�H��l�SPCx�Dvr�:����M�z��a2|��RE �B�7z����O4��|��!�e�,�o- R)`�Ug�H##>�(�Hk�p�f�$O�+�׳��b�?9��w�5��wa� �%g�\�?1"F���>N�`מ]��S�E��!v��ʨ�6"�8������4��?�Ku�R~Io�j��~!iP5X�4�4J�$ܬG�������iAF��m�\��Z=#��L�M�&�B����">�B�����{��X~Lα�6w27fjN���w���l,��	hN��X��gT�����\w<6��ێ�ۉ�r�-����/|�ݦѠY��\��r���s�
ٸV=�
�s��tGd��0�r]?4���^�{_�p���*qW�ut��>s��Q���

\�bґ�g��A��zX�#���`w�W~[	BF>?���H-�q��u�ep%�,	�mk=\D߾��w����j���,�i���u>�ێ�q�|0�����1�<f:T>((� 9��,0���%��h�q>f����mA�f
�|.���'��O�ξ,�IdɢDM��4������&1�=��p�/�>��פ���f��!ծ���Z�<^^eTY7l��dS�|NDn,�z�T�jj=��fC�����r캐���*�<��au�7b5LO�*ll7��+n>#a��qz@9�P�6��ѕ�IZ�Dˇ�P]�Pk;o���$�M�a�s}�����Se�'��[1;�l{rO|ê� 7��o�L��)q��U�s�R�ޖꕫ@���o'�c�>�fglk���t7p�@����DQz4g�Q�Y���{�`H��l�\mm&.�;r <tLV�L�N��X��-�̋48�Dfi�|��Z����r���ZС&�w$bH��ݎ  ��Ķ�V�D��{��Y%�9�:r�H�@�zFx��R�wZ.ow|�0�&ovx_߈�����y07�?;e�Z��m�vp�l1�{u#y[���S޸��#x�]�D�RkHL}��Mn�8_ �H�۵�q�X�+��}�ɳ/�c=�O�+�,Ե*`����9�)���	��Nh�N1+#-1�������u���e8�D�Ή���F����X�YW�eg�����~x����u�����m�L)Z�C��e�]� ;s���H	�)���N�L�z��E<�1����Fgƶ�+�d��l�c���K�	���Ky5bD4���ꖽ�k�=:���9!l@t�a�D,4�8^Wր�4�WW1�ls �Br*N4��h�[(���,R�.Z�ݐ|�*�+��3:����^�Q�N~(�*l��0~��ݑS鿣_6.����k��R!�ݓ��k�C"t˕�=̴�+���Wr�5�&�MZ��2�@H&�La�rG����&���<Κ��N��آ�z@�vI�B�_�4���fW&������N|!��e�e�|��Y�gc+��7�Ѿ���db�?����@,�(n�=���"��8A�H�a����w�;J����l�����YZ���j�k��ﾄ�FѢt�l��"Y�K��\�׍�J�bM󹍦띫�|�_���q!u�g�����e<�f��9�]7RɎ1Ar87�o�o�����"(v@�hR��̵���͞ǎ.��ľ�L�"At�4���`X�c$��m�	H2$I��S�D�@��$Z���ʶ�G��@{��k������_������^�Hu/o@��=0n���WX5m?����\����)#ߞ���p��HƑ��}�$���I���@/�����(��l�z�c�1��2cӸ����c��U�!�9��Og[��P*Y�n�p0�?:�w��1��3��SĈA.i�϶1�����<����_f���e�̲ꃂP�DBK]Vӗ| Fl?�U����<���Oy�a�
�`�"�u���qa��;�*:�������P�a�x�^@����^Yխ�Ɗ��e�)e}n�Qy�2�t����<���Q�k�Ս�wk�Cœ�.
m:m��Բqd�+e契��^~7����OW�oT�;�u�H�_̉b�ţ��zM�u��e8��aD@y0-��o3eݟ�,`�W��+�h��4@�@��5���7�[�r�i|߹,;���Ӟ���J^
��E���f�wV����F	z�j��6Hdv�M"K�(���sX��R�W1�zJ�ԙ�{�lZ��5M��5��t��۷'2���G�ry�?e9�8�!��t�Z�#=� �o��[�3Ŀ
P���X˝ ��	��a�P��@���<�ꌀ(Je$�;�9F6PT����r�c��r6���Q������\� ���3�NmO��*��4ϖm-&�i������w6�`�ɛ�"���X3�ط���
�m�m������Jƪ)���X|�M���/̷`3�I�\������n;>�����=��nnG=-�í8�ܮT��͗����|��S����Ɩ?eQ�Ҹ"Օ���Α�A�Tzԭ��r�W���1��1�C^j��7dO�}�2�����������f�<V�W��:�)�Z!�]���to��|S�AZ�k���y�,����B�n�X`�q��s7�i��/���@���'FT�˟kc1L��E�����1Ѧ�k�7����p��X�w����tgA�AL�c�����s���1 ]���	]���D��=�A����A�3��Cm�.�Z�':шɑR�Ym���r�\<�Hr?������s�̺֐��bd�����͎�sm���¡CI���"��Z�Z�M�-G�Ir��	Y�G�� ����G�[��e죑*�Q�8��d�J:��r��')�ǅ�~d2o}_�}��Gzh�v��t�(ܧ�W�Α�&���Ѵ�0"��K|�Gi�aJ�����?�C�b�p�����/���2��Z0�Vb�,Zƹ:Ӌ�Й⟩�K2�	�X�#5{��q����������v���h��l�OǇ�W�TA�~K5X�ʝ��p��0ͮ�ɝJ�ʆ��.񒙾v��^�D����&˖�Rm��+�f��qčPN3����0l��׋; ��m���
�%�e�.�(�jᓎ��`��S�~�X��_�ԝ�����[<���w����7�`��@�{w7=��=�V�⏪���������Ѫ�DEJqnӴʘ�0���EXG�jIq�׆O�������W3����$a�Z*<׶����t�&�+`����<�(��Z�ҚN�L��{��|Y�K�3m�����oY��B�Խ�+ؤ<If�-7��-q�?6ҩast�F�Zi��/xk�;�ex��{5�ʊ�JQD��#�<��$�OP�_0$�帆��]��I��$e����n^}��l����$�f��I״M񎙵��L_o�y��o���A�A�l4��)�-�Q檧t����?���E�l=���w��pk��۞=�����|K�P��o���t���<e�Տ��F�K���Qf�����qAP���f����h���V:`s\�]��O)S ��_�mE�7n�#�f�w��ɓ;�>�O�d�.�(56v��ȕ������x=�%-Ȳ_�	��4fY`.��Y|�q��"T�������k(���4�P��6u?*nBL�E/IX	Y�}���|{)����C�Ѱ宑��<��X�A2Ej�f���� v˪}=�����!�?}9{�L�!5-+~�g������'�c�>���u��6�цD(�x]@�����b`D���q�g�>C�Yx�\"f�c*��.ξ�Vi��`O��C�7��q�����`��SW��5n
��Ƨ�c�J��gM���wk/�S~06&8�_�~������!�(���m�R6(B%�
UyMzc%��ƂT�������״NXN!b�|�qH�Q���0N��=+[�S�&|77OQ��6O�̇�3ƽ�9����5Nm����즾���L��X�fy�5O+�����M�$^Zէ����K�� T��{�}@A`��n�)������>�茶��8l��)�����m���R���&^�O���H�N�x��@�md*��g�E)�6f"ĪV��ט�z�6�'h��T�MOwql��1�h$~�ŕ���9��]������V�i��M4r1����׸C���%�q)��
��e�v���1����>V���+��ʡ-��c��h��6���	�Gf7��(��͂Cc�	����jA�������M�1�?�,@h��~�hc���q�]�(O��e�ԅQߝp	���r ��h	�}s&׸G�m�?Fa^5H��'�Q@�q�0n�Ϸ��!{���W��b�l]_�v��Dz��<��������ǋS�4�w�:�!�P�V���|cP�]�,�	��񕋈�G!:\$�|l�bY��Ly�l-��
 t�X�1\��=4�3��a�N�j)��\�OQ77��y���=c׏'3�nDf�Ï���Z�<¨�Ŭ�u�G'�A�M,	&�����}2��:��e9?���(e����7q��/j7AzTN1���֞nz�{*i|�-y�S�K%��:���K�ǚ�|o��a�I��Z������Կ�`��Ţ{��\k&e�Tw
�ݩp�-���%�B�k����i�JC�-#���UV��X7���b�WW�e�x���\���#�;��k�j��f�z_T���|LD�a<2a��W=��dxb��gmĂ�H��
ŋe�`Mm�kʓa�?e����`���-S����}���=�=n�9���+�
�����.�a)n��ӺB�"ͨP,Ġ�Ș��������M|�{E�op�
|�|���Y哽&�PD�WV�@_��ot�Թ�����{#��r�DR���I�D�3�2��/W�/���ķ[2�;�}l�2�ǤV!̓`q�+V�.��ݜ��y3����)Um@�L����E����W�*�߫��;G�;%��K�X� ���;�%c�5j�����2��N��y�^��a:�ta���G��C��P[Ri�0YWt_����e����R�� ����LC�T!��7�Ӧ�|���l�O��k˕������t��/�`����L'�Oߣ���/�/����|�@�u|x�u���9Vn�>:��P�^���f�R�b3�������kvz�P_u5���ӶRf����O.�R��W,A>{y�Ə���Ñ$V����w�N�6'�\�GI�T/�g��0;���ɵ�f��~�52��T���iF|Ð�|A�-���)�x�u��Rn۠�U܌r/&�D��f������;zwmG��N�&����m4��9���o��\u��m�SR0�҈�J�֦ ~\?FE�36�\p]�EqɆ/����3�˓��b�93��/��C})U��� �7�ɤva�tC��bsv��k�`���oR�YR���S[�/K|hW�+c�`����S4����-�34���I�\p��;�4χ�$QN*nԣ*�/f�,T�9��d~����D�kQ�FpB�[=����$ʺ(�D���1�@&؁I�Q˂�V/HIi���>#Pd;�2� ��`��ұ�k�*����:��Ѽ1x�����.V#�l����*P�ݴ{�od�ѐ�t��3�7��|*X��D�BO���]9�e ��u� �}w�z7�ͽ������j��C�����ju?�;��)���T,�������t���o��)7�����7�1���M�9=����Zf8m��ڇ��K�!���B��)4 zӱ�։�0�>�y_�U�o���cʬ"��J��9hdG%�1��\"�3sUĘ,�WQ�t~���z5<=Un�*�b��ٴ���xq"C)��x/��y�yR޷Nqz��j��MC�o�-G�=`;�杰�x��/�V|�+���7��g7֎{�C���Lg�w�[0O����Lʇ�H�t0���v�_䌩��NU(0]Y9Кe>Ke�^�T|����>�<�|����}���=u �;����ة	��ϼ�4�<��l�{%eBr�)�PS�� -x'�M��lX�2,�vV�~��M��d'ɥv��o�3����Wa��S",J����v4��>�G��G�54
�!�c���i�H�@n�ܯ��b�b�>aб�X��$�T��(��q똑��&���� Kݛp-��]C���i#�[]9H5��ڿ���˴�&8Q�U����6z��o���ǥ��>
$]�0�;O��O��1< eZ!~H��֪�oӮ�Qa�M�.�r��CxA�S+{���7��^����Y�!�{M�� �4Agb�'#g5fnu�,��݁��҉Q��B����2$ɂ��2�d�xDls�d縚���a���ߣ1�鲹��i���-��VS�
�b[\ވ�FǬ�RYnQ�o���C���wUk��*�v����:
��)��,v}��g�jx���	Y�N����7������p�����1G��QZ2��п���}_3c���s��������W�s���E	�U����]�ߧP�S�:��bJQ�#o�F O!����ilg���������#�2�1UP�&t�U���!���#N�^�u�Ԗ@	�h	��q��M�,:;bdCX
����A�?粜�}��Z���@8�=�V�*��tS�t ҋfy9�`ӛR)�Ѝ����U3�7�G��ۋT�\�5ѯ�k��|�']�\�S
�����2T�G��E�
 ���u�v@�g�����>�����>�_B
|�~Ǣe1����4�^�$���w�4� ��Ic���$��k{}������n?ϝ;�\dDm)R0�鴓�$�V����ODw���F=�(0�>nb�G��C��ʣiJKR�yLY�7��{J��` ��⋎_ݾ_��{w�a�:�̐�萮������Q��U��U�ø����\\|�#0yeo��)����?|Q~�*S�eA�Z�Ɣ�����]�q��ҧP�^#菇�BjHՈ�Ng�|�ev�Le���;\bב'~��� *�������þ�AdZ���8f0�#��|�~��A \! kXkߺ�pnP��!����hy:,��ɞ����$&j�t8S�Yh����b#���-��aM����]/��E�������a8���lX8o�� `|t�1�Ql�����O���S���E�ݩ&�}��&#���5��n�; :�޴/�h�W�@���X��`<ʇ�TNh��o�
����؞u8���u��jܶn�cg�������d�i��_���}P}��������muģ{�&�~����@����jS��<������[�;��MOC��VX��V	���@�8#�JZ`ض���W��2����78���F��KA�فn��[�g��\��E���r�xt)7r�Ie1��t+A��~Hv��� \����7��p��x���[i]��L�4%����(*}����g홗���[��lh�)�}�[ȝ���o��9	��]oU��l
�����L��5��+S��t�o�]�wSM4L`3ngDt@�av_�@o��,ގP+����y1�=�;�MŜ�N���ֶ(~�d�p� ��b�Jla�ŷ�e��e�NX��
�� L��;���lyFYob��-X}g5Bn<ߐCc.��b�µ����$h�����~RlF��'�e.E���U�^�]S:R�_�|O$V�'��_�1����'b �~L��?�8\�Q	p�慄��bB�5ARJ����T����G�yTfL
`ZA,��96^u��}1�1kM�=���_w�3@4�q���3-і<ʯ�1ږw/ 0Ϋ|�q�GEVn�ְ����;nT�i��ړ�����	�L����Q�Ȑv��_�{õ���'د(�l0H����U"�z���d �+����AV��dT7�<?�'��îuiX�}4�{��H�}s3՗ߌ����l�v=Nz�mH�z�-ׂ�gd�0���ϯW����1�խ����sS+�I��-�ً^��.�FPS����Ꮘ��WI��PVk^s^Z��	/vƹ�q�kH!�8�%���s?�.�˷؉5�P.�s��Tn9���A��!���N���S�Oȃ����YRk���+MH[��C�ťx��(��g���n~Lz�eJw��AS�?�,�b�U�Q1����RE�> ��G�e������?FB��V�m]P���4����	Pcߡ�T����*b���h56ikZ-G���{�x��fX0c�(�1:D�up�\�÷gٺ9�8 �����"�<��R�F����E����e1\T�ٽ�f'Pӯ��I�Z��:�,ٸYN���:^/-���ݯҜ	g�0{�)$���w�G�
�m�e`2��L����-��DӄOhJ[:����?΀v���v��={/���}��B�P�MVq@P%�]��ei��[I-�@�a!���Q��pj.�\I�h8M����V�~h!H{����xB�@����	l���Jw�c�If�2�	|�������̋.���lC�.%$�7�:���ChBPxN` |��qɜ�0J��ٮK>�t����c�噅�j�?j��!��F0)WOR��$��6H���|o+a�����h����M`�������K#�"��Q���RA��F6O��D^&�c{��k��u���#��Dq9�2o7�Eu�c��	#��}@��P+L�D�/��[����Ү� p��}O�#�kFc{����9�����Â�i�,5�8���n<6� G�?�P9������t�˭�k�#	��Ii��{�M���C�ь�(��.�Տ��LCn�`"����Q��b$MV��	��	�_�g������<>���G�uwwA<v�SE&�#��1����B�JV�mS�q񊦗�%��p�빌�t]\&�����zb���B��9��AoPc�Yqu�&��o��nH y�� "��H�Z��t��
͓xE��;�9(�0O��s�zv����]�32�d��+�ꗖ�U;.L��ڮ� �A�[z��h�ϖc�9����@�i[�aGI��o04�ø�dl�HRt��r�İ��ic�7e��TwΐBI�X~�`�g�c����]�c�L�8�XDE�6�/-Us�hF�^\�͠V��
�������lQ#|�(,TZ�酯x3�`I�&-��<=ur�3q��7(��>�[�����dA^(���(֎q�;�Ms�p��併�D�p��M�%��5i�/��6q-���kg�����1ĉ����"��I+���
#�0f��be����X_5t���ұ��t٫Q!��.K�a�Fx��3��f�������k��)�-�R�K"���%��'�v���Pl+8�l�<(�!�P�,��]dǲCM�N�ڟ��nk
�����l'�ϓ��OO�{:h
 Mgk;���� �3*&���P�d}q�:��@��4�(�Ò�tp�) U?�Ҙ��4��CFoƶe��W��El�e�!^Gk���K�x�j�㧖p�����;)N�G�2���w�����|}�ٽ�� OE\��k�a-�p��-���f�������v=�.iz/�2	iH}8\��M���&h�����8��Fq<J�}-J�ǅ4�:�jނ�x,��۪3���ATj?Wl��,���]�3������<q�#{�zW�l���{�4ޑ�� ���Y�8�VV���O����{��/��^�>�wvȊ�md'^�g����JTVa}�`�0�)����tct6�SQ��iԖ��+ �5��;�_~ݱR~��0G��^�bd�]�(Fh,�&x?�)�~6��ib�ɕΚ8���k��2nɦ?#5cT3���Rw�mGn��&㨬���t�lzsV&m5�����1��{�8y6(�6���Y.+j�`�1�\�.���������g�M���٢?#Y��������#����2�_pE�$$�Z��g�z�6LM�y��c�C��޾i�
L��6�F[�;)�X�ųx����.t�g� ,��,��cf4�T^�G�7��i&4#M��I�T�pҳW(rݎ��vG�����O���2@>x���?E���
�KZ�1nb��ѻ,,�pSgj-�Q����b�;t$C��@YH ���{ɿ���0࿰��-&���|�8�h��!*�#M��C�����"o�Ts��̡
G6��PqQ�����.�0E��{����&z�/�Ƀ���;+y{����q�-q�6@I)�o���MA��E�_vu�9V�Ɍ-"K�<�r1���H��WГh*�O6l*�hZ�����is���V�K����٘�;�S�
c�&OYA���<����M[^*>|�1������9}�^��w��Jm���=�j��uN�<H��B�X$O�A��h�A�8��L+��N�å9i�a�H�m�z!��F\�< U�OZ�|z��ݍ3����&8}y`��5	��Z��N��m��.O��'��v�d	�h掽o����򎅺u�K
H��U����@�T��X rn���Z�`�+E�+����v�(S͓,^�'�ƈ@����4��_
��:���j��4�D�=Wg��G�H���1(r��<���i~�r����}�ʴ�A#R�B�Ȣ\r��e#p�xj���r3��zao?o�Ϳ�ؙ?j_ֵ�OFtXs���`o��t�'���[g�-fN���ݝ����A��N�v쭅7�4����D�����GL�÷����Q;u����ӂBG��k];�踮'#�j��~��2���gT����������WF��^M������:�v�ޏ& ~PK)c*	I�u�q{�e���)mL��p�	��E;2����O�0����HFY�x��O�֌f��~�P(<���ܸ�(9���� s�_	/s���M���ݚ�V$x�1.��^�qJn�AL:f$:�u��ǢN�k�s�ui�
� �m�����%WE�/�㲄�����Y	�P���d�&�pΓR6�����)c�2��a���( "T��N<�|mP�t����P	+��.���,�����wL� �W6A�}@��Bh�P驳�wv�A�UV��e5��}�ͯ�>|�������r�r.���z3�yT�/`X3M�JH{����Z�����ѐ����Ѝ�b�I�:��7�ߎ��;�Rx9�o�G�j�Y��,���'�E�HKCkxY�E$\��џi�G���Lє&;cX�h�G$��S�u�ǟt��Q��&�U8�i1����H�ʹ�ǻ�\�8Ѱ(��g	KZ���,|�4K��m:��W�|]m!���[q������G{����k 7΀b���z���t|��4[����#��g�j��{��?������{�A��tR�\~�n�������)��� �U�F�jo��*cq�ѣv�m��P��������]#�j$S�^�`�±C$4�,P�
�����AN�2�Fp�a����ʐ�|��I�lJ����)����Ćl�|���lH���b� �5�%�g��L���
��-�,kwM�f�.�l�sc<8"G�>����b�6���p��T�'J��>�8}5�x�)�1�Ku�^�a��7�WI��|�ġ_����ތH�98sJ�)��[jA�{�)'��&�6��2@[�<���/dBoq�a��!�hx�-��|��7�~N�K���\i����>U;>�Y���$���Uw!���m���}�T&��,�Ap�49e>�"_����ں)U���O�؄X�zp<W��3m�9����]<�|z����=zv�檉�C��-3*f��1Q��?�ROx�G�q�֤n5�>�w��)��,����ל|�|�+�-v�ʖ�ޢ��H�\�C���M
e�p��"X�� ���Y�b���/�����>��~���9L���pa���d����:6�zx�9Qtq��cv⣟��WE_h�&Rf�����Ւ��m��3��{������,�`gn0���I��N�H�C�V�:-R�/�]��vbuh�|��%�i]��� ��Co�'���-س�r�Y�,ѿ�f��&\䦇���Yy/�ŧWVy(��z0���B�XsL�x�_��6V�ѳ�x3Vu�^:��d3U.�����m��!̑K�����?tIw��uz��6�X{�V���ƈ��;�ҭ��5j�v_w�X����V��tS�fZ)�^��1��,�^/�(<�^�ڎ�|�����F�Ռ�%�ꕲ�-P���+XUѸ}0T"K�e칱�K���q�n���с��RD�1��.%}�)��K:M����YpG����FK�����e�N�<&!�]�s�_ҵ�����Բp.�}z�bH/���aݢ����s8��<��7ޭ�yjt}�Hc������6�pG{;��ث��t�-$�~�~h�|�B�	|���fT�l [�a��Ϡ���B�Q5�G�B���x�׭��g�/��|�Z��v-���E�)J�^�̦�/N#���}�HF�tN���c�Wh$v����oa-�������E�nĺH�A���<�<�s�$A�j}�H�FRl�WX�˦���n)�0���ee�+B=]�c�8hSؽ�R�l�N1�$������u���N	A�;&���o��*�i~�2��݀r	�to-`�AF`K;�e�^PA����'����.k{\~�1�g��1�p"��U��0��!Q���T�к�x%��Q�&ה�����2�8���z�MvY�푨b�Ӯ)�٣T������� �7nZ)BH=)�2����c��M m�A��%o{W�ͯQ5��nUM����?4�� w0��
�I�tS>�N꫒��K%����F��A�l-�)<�V�ܐ�Q�3v��uR59���z�k\$>�(	Ϋ�~ͽ�6+��|�?�*qٕx�w7p񫖗`a�5 \� �9�2�%y[o%���s���D:ڿJ� ~�X�z�S�d�ҿð�Ќ�g�7|����'Qbįn�9��PR0b�}�Ea&B�}߂���ѩ�;u��Z�̔�7�p�<٧�`��I//�_�~v�F`�oQJ����화@3F�������!Bl/�Oe�,��۷��1~6�� �� "�<?�-Gu]\ �ގ8���U��̷a�A��f��X��%v�k�Ҿ�~CeN`XT��z�1�ZxE*�BD�y73��iځ�Ѭe�=���U��x�W�`�g��7�nWH�=���=����U��J��r�He&rϦ����ޢ�)�lX�¤��oIwl}��+G���5�L����G"�>>rm(b�2�&!-�u+Sb4QG��,��#^)j��M�_���Gb�z��F.�R����2�A1o+s-�?$������=��5�&�b5[�� �olѣ��]mT�	�0~�D��J���ߔ�ofKߩ����WΏ�ϲ�j�2Vo�/s�Ƶ�82s�)!4o{�J�|d~��S�Eq��Z��$�!|�Ŷ����Y�5�1�ts���R���.,���'��o�8�,�}�e߀B��"����V���#t έW��a���e���kB���R�I�uˍ��c�EA_��r�!=,�5�Dl!�E<���Q��ҧ�[�82fb����8�a�t�~Z����L��tw��DO��A�ed<��)mҭR���~n�g�"#�[�'�b�e�P�h	���Z �a��d���+}�Nn�h6e��ixʌ/)�U��m{FվMIȨ�^�>}����j^�	����(�M��_�d��������w�?�'v*;E�Qo�=i���-�Y����"3�	b}�.�=3�ȩR4��E��\Aô���N��^�/��R��D,F�o�~�;�MrN+�O���Ӑ�I��V�Q��[L)+p�l	�1�O_�	�u|��4@#��`�W�iQy#<'����^��/����+>�⢒����T1l6?%[L���aXP��pԷ!�s����.$�
���&#$��!��f���T����
�,�!R�o�Td�Հ*����Npx�5����s4ۡ��C�50���"�ޣ���Ŭ�oB��-����}%�)������b*k|�14@�e.Ԝ�w}
Q�I�A�qջ�I�Y�x9��o||p�]�1��tx�?U8�7Ia�VɄ��!���	K0�V{�p�.hLԀ:s�Dc�],��
�};{��]�Y�ԉ��l������c%���LI�RI��O.pN�?����lj	o��M�/� q`ᮼ!Dr�����ƴw�w��=�s;��p�mv1�����֢J�t��"�D�V�z�R����i�����㚂NV��
�s�OAU9}�!����QY��~7�3D�zB�HA����^�b� �~�%"�V�0�0U�4��Mc�E�a�_=4�3wzR����2��߰��V�!p(�ǳ�¾0B�Ds��xB]xrI��ɕ�����kb4�k(����.����'�O�<Q6�'s��SƛN�.���H�F��a�9��AzR��D���6wn���7���2l}�Qs�ap!J�@P��S������R�y�+�u���D�g��K�u��
'+�ӆ@I�lȰg>{jZ~d�������d��3_ڻ*Tn�A�0z�y�;�w�r��ux���m�5�C��h��u3���y}xy|� �Iz�3�n ����G:�9 n1'��M	���<�rzT�D�f�,*z?�`UY��P�ۇqS�;W-oJ���|�s_�Q������ڪvqI�~�νMa��*�3�&�B�b�Lx*5����:��"�S�=�	I�B��a(�,���e �事�����]���q���ʀ��*�	S7R߮C�C��"�d���χȔ���[��^���U��s��b4~�3��1��j��@p��}��~pH�_����.�)�����$�6/�Ɗ���4FB6�Ns��&C`�ӱ釐B��c�PԌڨ.�R��'}�Z��Ã &O¾�m���|g~c�4�H��O\��K�F�f�fӏݗƂ��1V#�_�N�5C�y�{tD0�t,ˀ�77/j���� "U�ݒa���*�\>Qͅ���ƍ��{�ֈʿ��$j���	�_�_$��{A=v�R���?]�&Us*{��o�� y�����oߡ�$P(.u��NQ)��kG�W�#]� �p6w4Mc�<��[M�ѓhK����d�
�N��S�y������m�4��'�]�3SFM��Y{�T�ܳm(q�h��^�|"�
w�y�A�믿cj�}�Ҷq��hԌUg��Q�8Qc�{S��*j���#��7ZWU��K<�B����]�l�j&H�E�x��hK��<�h����-R�����#��\�p�-y��y�X��64����b��&|�M�u��
dӃ�Bg��$�D��c�(�b���㌭~�����F=�^Ԟp@����V�"w��֡���v�k��+I��̫�,�  E��=	�Q1��Gz<�����`q���+J�'�Ȥ>���v����!��5��/����7�"Iѯ���p�+���q,�o�n�6d�rhg�1��=�+x](gin7�qa,�E=�j�/�����;f�J� g�)�?4�d��0�N�hgQ`U.T$��<���p���Λ�Pͧ&��֊�y�z��H$y��:��g��i��iD_�b���^��؁[��*ç�����)��!V3Dqҳ]�U#c�8]��i��ea���rh0jl�{4I����M�ܮ�Kþ䕤>C0�����v�둪�h����0hUo!��o׷���{ٵ�sἷ��v��-�fM���o.�Db+[�/�|r�3奛�"��[&�����e�m�9,!�%S��|���I�W�9�k��A�ӣhBT�_-,��)���?R���&��	b �vL��������n.�G��0#�F�l|,��+hz��vi��"`$�d��!U��J5�P��ytV��q*�;*�!�py�Q;��;������R��k�r���x��N�ƀl�sv'��ѭ�'K�.�&�=�C�WY�.��#�-�#��U�����e;�A�r1B���tH�s,}�˂H��/XB���m�����~f�^��R���O�},F�u0Q��Y�r�aU-7"�"'��v�Oʙ�i����k�	���B�x.���V�Ro-��w��Ч���4��\Qb��]���}�|q���������iiZ�'�r�@S��S����6�_#�am�fl �Kb�3�%N��U�}=;P��~���eҲkBEj4�Z�,<�����!pA�H>��ft����r��K�޵��.yM�/�\:�o�"i�a�@��{:���2���ή�Ʈ@O�F����L9���B�(�iK�M��u�X£V�X���Sj"Y�n��9G R����6�gپ��g�n�U����k����M��{�K��D�R�e}�@�7�aƆv!Ih��L`o�+�sϻAc�oaX�����K9�����ot$���pebNb^�h�e�ژ>4+�F=sA�c�vN�ϊ���� �0��]
<�B�y�2SK'� 3�@��K��OWd��V�0��2�KrS$�Q�p�	Ā��Q%θ:�7CJ��j�0E�g������������.����ʢe���:�'D
��8<K�@$���Ɠe��O�ʮSpȍ �./|�V���I�'�c9~'�E����Sπ�i��}1*l�(��Z$�aE<:X����[�nΪ��z��{���%����Ҡ,@��ds_Ƚ��˖��OX�XJF�P�P�F������jt�\�Ҏ� oF� k���RpD�`���β�,��Vz4|�����2��=n��5�U�
�'�y��.����G�	��?�pp����¬���=�jl�;�L�� �}#�G��0&��1��z)-:%}$0��Z�,�SA�I��mk8�N����&6�~[�,)ȸ��1��H�F�X����(J����%���DPz��,⨹N���zj�Wsx�!�

>UH��#c8�n�0^[;����;G"�Ү �-'�I1�����#��YR:6�C:snvå�=T!�Gh��_�K����)ɰ��TD>wԥ�!�}�
ؼpU�MKE�L7>g��<:Q������t������y쉎���݀k�ǡy��
ַ%�}_9ˋ90�y��5�Oz�m�b���y;Al�����U��Т���qJ��@ٓ@ݤ�����Ծ������0�)��I��[��'���w��6���x�n�#����%�%�	W��>�Ԟj���}n4�39;Z��W
k<��Z!_���i��n�1��W�2���4�6s(��Z].�d�9�0����j���sA�)FnHi���nW����%p	�*^Y&4��T�A�6X*YQ,�ڻ�Fe4�����I57�:�5.��6�Lf��k81�
��r�+9?<c��P�2��l��w�z�q^��u>��Q�Ѩ�ճ	�N�\p�|�p�md07�ځP���k����|�F���%�F�7bК@J�,!)o��G�����~-��B���@FNb��q7a��|Tr �RVͮQh�������t��1�psV�ۛ��q��;�F%�vXu��WK��#W�V��E��,s5�O�ů�&K�|�P��э��`Z�!\>i�c�&���h��3:$�)�l[؁E(\�2Д�"h�:��^�%NÊ���+��^����jX�m�ۅ�����UPT�O�����Bv뻵�����j��acN�"�6�jJq�g�2r�0%�a�6t��E/-�ԕ^��[ָ�cs9�z�UsWb�� �'vJp�9��N�&�����t�d�"�0�Dzf)*}���B]� 4G�rB�rkt�Rc�р�U��/gn�Pp�h�,�����k�-=���0��y(�|vU�f'�F+�ry��oK`�����0of��tu*��M���e����<ʻ&��6�)Q�Y�"�+d��g!�܏ze�E� �k��^/Pb�+����<(���:d��P4������V�s��,�4K0����u�y+�Σ�V:�ې��K���'�< ���it���Q���~i�/rQ�m���^�W��B��Ǘ� 9&1Y�Կ|3m�O���fVd�X��=|���N!��.�J�$��?���x���Wc��p:�)��Gg�� �}{îӮ#u�h\W/��YG��G���fC>5�W"j9)o�Q,>�
1�����d�(�44�c��ɧtY��.**4y
kjO4V�o/e�A�1��@ �5&ҏ�h4�EͷMz{�m�F0��K/�Z�m��E�"��陁0�j�>P����a�iG�utY�����F ��6���R�x�_1�^c���v-�<��e���	��#�T!Pry�Y[��ˁ�퇣��4:m��8R?�cS�g� �6�R��e�<�e��1�2y`��tb� �ϳ�����X*J&".4!D��x�Nւv��g�7���K�	&�E�tlK�x�a,�h�w��RTONo���l���V��7�q�$i�09��P"�^�$��ٞ�#�5�n���zc��kV��<�-|�v�Y�P���/=� .�eHC3���ʸa�0���L�ҏ���IG(k��@F^��a�2���HP���R�]��huP�-	⠶�|	m^HY�*$�y-��'��Q.肬)Q�dSsU6�E0E	�A%��T���P�����썌2�O���h>���68�G�0y�,!Lf��'�E�`��w�Z���(;�j��8�g����P�{N����XX=�e�cq����w�ހ�k�iu,�!���'�'�e�J΃p*,ָ�!���_��}�	�D���Ex��^@�O���[s��jY�v�	�ϋ�qo_",�*W�"0,;+;�]��b(٠�BSp�'��-A��R����R��_�����Y��ꚛ���@4��_�,E���	��F�V�vX]|�=��#`�&4h<ܐ�g�ɶ�s�tl���T�+-� l/tb4,����54#�E6����Ȧ��$��4��%��M�-Bʈ�㈥��ɦu��fv�q����s?ng�6]&_A���pU��(���2ڕ�C<8ʃ�����AV�<�M.W���e+�QL59�z���}$+�وFsX����>� A�0������l\��dG��ⴏ�vGBA����3��5�S�z�I��M9 ���gZ>��&�w�l��]B��w]����r>u0%
M�!B'���#է]�7���BI���U}:�[�N�i!)��g�b�� q��R4��'�E�����W��&!� X#�Dr���$���A��[����:�,��-��R�����VF�Lw����¯{��P���H �κ=�����%f�=&Z��A�{֜�W����p�v&����pc����0IX��s��l�ߚ����S��'�Ea�a��$�yh7m����]�>	�#�ZhE�C�W�!N}�Ԑ�r"��ȓx-��^hB� y�|g%����(u�>�����^3^����7\���e��A��[�!_�=�.�fnKx�J����*��Ak��ƣ����4.&��_!�2�����K>��V=�m7ߞ��P\��hE�F��P=���z�s�A8S�ޙ�6�!1�%�k�$2����@&ﻠa�@V�X���v4n6D@d�_g��"�N(�  �G��Hg�d~�Ʒ�������#��t���6�����������x�8Bz�]5�E�Z��@AP3s0��{�W$!hP�0+�����p��9V7� �����!�n�\�w��#m+�F4V���nLdhdC]#<[���~��ed�FV��W�r��aD�����oB/Y|=�LF�,����[Z���I9��'�4�{��C��5O�۪�B�|t�C��	�r��/�1s1i�ĸ Ó���n�����䠱L��x�B�?÷�sʮ{�h��ZĊMGk�RP*I8į0�� _����{��1�Ez�AU��␻��>�����B3-�bP��]^�V��0��"�QpـaU��"!��*�����C�KBa�BO>��{i�\ಬ�oJ�� z_n�~�QU����?�L�~������XZ�:۳��)�`�N`3��%�sn�1���$j�^Q�B/��!C���W�HN�0���EXt�Vݟ�6.��p��2QwL����*��D�S�ʾ-�XA�f��	�ks������C����n����!��B|��I&�X%���13k1I��U�ѴU�%�X����D �W��c��§a�5MUq� lE;G_ɃU���b�!�=UЗ����շ�
���
����K#z��tD���/9M��B�(��at��c��k��u[Z���@*3T�D �܁Q3�bX�z�߫���x�lu ����-(OM��/C��Y�A�����{���fh	vCrU	a��AA�%!"}y�g��=��+/��A�<�͐^��K������X�C� >�8�4D�tB����Ok���Lw�E䱷��xM�1�a<�d����QPߊm����.ϤMf��&# �8K!y�����P���i�|����R��p���f��ݮ%�O:���w�c�}������n9�p9e\�����j��@��^i������%W��j539:h��T�k����>�)�v�Y#��sK�I)�)�f��W��}7� ����m������I��fWf���|���@�"D.Zto &��9��eI�C�M���5���Ó�'�]�I��J���sNw[/���e�Cp��=�h�:�;��D�,����~b�e�!v���<Ƞm@͞�X��dP�K����=7_�lqG��b��:�=8�&w���H7�|nh'nH@4�-3?�'ca�-*4���լ��$v�u.k�=�K+9�n�p1��?x?�}f���i	D�*�{�xl�3�Ik�ć{�p8F���ΤÁ�Ła�"6�G ��*6�S-�3�;����"f@� ��Jz�U�Z˫_ڴ~�a�>� Aa� ��G��4�+a��Q�#A��Pa8�k߭&�n�dK�}d��-�h^/.�s7�p���ց�_~��<0��.���a�4������uQ�ܔ6�Vpx��ADww�σ.��3�:��Rs�\XS����?�n㩃Z���� ��ЎHraND���#>N�F[��&���Q�`-z���8�#i<���e�B�,}@~��Q�(^�1<�y����:��1�VV�� �]��bl)Nc�']-�#�r�5������k,�XL�u���6�<�R������/ҊP5c��MĖ�Q;��ԥ��-$[�@ �@3l�)]6}��ѥK`�jp����aP%�%�_��m��P~W��Ht�,����~헋x}T����3l�v}ԟ�'c?s��	&4�C�,��[2�a��M��e���	���/� �/*��®��N�����?�*��.�ዦi�b�`8�@��9�$FG���1d�VȾ%6��t�N)��_0,���u�[�7�<h���֪e�[��gZ��0�����������[9�
�|�������s���Qe�H1�4�促 GC�6�O��
�b&�]n�����^�!�k�K/���N���	��8q��9��0p�~��|�vY��'Hi.�����ZWk���"����:�Jwhnl��������t܋Q״�׺�L�C�̜��/�;���������B����v�e���� m�h�.+ǒ���p�"�c��6��\x��Af�ا���!��z��:u>E�x�bڇ�zA�����o�k�a�����)]��$n1N4���Њ���*�NCO&�7m.�y��z�rQ�;�B&d��pH$B���s�I���w�<�$~��<�Y��@���&«HX{٪�6 �8f���ɨ�C�P//
���Fմ��2�b�UQ�;�G�����5$J�q>��"~�<N��f�t;�L�پG�b��#-h8�_�K���uPK��],�[�3x�)} Ҹծ��Pz(�f5���()ڡ����}l���~��|74gY���S��)<�c�j/�
kv�B��=�-���Gu��4>�=�k@�,/��L5ɟ�l�];}0���;�E]nF�粿���0/�nŞ�t3�x`�و������E��R� `��u�\�.3MC:���9�2̦�>s]�xO����y�S�(QQ`K�N��>�S��b/4T�yD��p)H^�S���m[.��&1ny��#-���\������U�8�:ʘ]�`�������8�c�?�_�O$���e��>��%�DevE g�֔d�L�Ry
�$?�1p���/uȁ�W/ �]O�{e��P	p�-�Z__�5�k��P`�sd����	NtJ������2�7>��\(J()���>�9�ህ��ڻG�=�*�L��9��v	�/�tx��)��B\bs<�e�5��L�� ]�}1��.�%/>�ȳ;����!*�w��-�J,���<g�Y�<G���=f�̏ 7�:$�k~�}$��W�n0>;�X!@J�TZ�P��������e{�z�sb��9������y$#��"�!W�!�g�25��gK�S��o�xR3PI���]y�$j��y>l:�K�m�k����f��5��ef�:j#R��ɗ��5w��J�� ��X�^'{|�FZɦ��G���8����LϹ�ޚ�IK��#�U忆��d�p�}NqŮ�粣��e:0B�MX'�<2W��Q���� DIb���D�oi�}i%�uH�DU���`�q��Y��+^����M<~��|"v��hcն�ʉ�OTC��`�̵�����⏾��I�c�n��\�
�t���U,��n)CvF�0
gRpO��(�-X!�wf������Y���+��m�_�b�v
�:_�Ҭ��7`@�|h�@G �PtK)�"|������Z�yLX�EqF��}8ڣ#*7������r/L�es��o�Η�U H	+D�6�rwwLk��Z�Z��jj[���p�gy���4���ԯ�C�V0����6r9Ԉ`q�?��WImx`�;�f�VV��j��JZYl��5V���H��˗���%sU��"��j�_?)����-�:8��L��L�e�LǍ�v.�{�����*��t���~ܔ�%�Wr�N)����#�&(#!���:��@���ᇀ�ݭ6O�IQq�d��~������3ݶ\��2O�j��^>��Ȥ���U���8��k��4�n-�� �s0�)d�6�|{���r5.V�Ɔ9���X����\B/u B�_8�
���^k���y�B��t
��{��]�#��سM�`,6�Vh[��"�j;6SO��uI����*]������r���l��ls V
�o�#O��*7�r2��B*�k9�ѿ�r-�2^_Փ�]���z���{ƩMZ�ct��3=��$��z	��3��,ը�k�E,��qoAv�A6e�ଘ����c4z��у� �(��'3�)�誱ii	��6'Ha���ءPv]�wv�ĉ��S���TAxM��:.+���U��h�<H���ˑKa�M3%m^�wS��ݪ���eBAf��<���=���-��Zl�kI81h�<NM�S�;:H���+K�O�YG1��c��.Uc��͋K���6�������݋ v�lN��!�qYf�J&�H�F�sz>���0�B����E��U��V�7�}��Z�!≪%M�a��ԫ�,h8��zT�1pk�B�5'NT�����"�B{\��qKI�f�n����T\���xߚU��|���)w�౵5A��Bф�~��BI2�Z�ey
�t��R`�dꐐ�'&�X����7¤���l`v��Y�>�?'MSKr�헽�N:[��+�	د9)�1��㟷��+�B�����ow���P�\/�[�4"C]��\�АͽM��2 p<�"�1o>T�l7e=��{��+vI0"x�Iw������>�:��L,#�v/�c����P��<њE#��_å�%�Hkh�@B �8:\F�3��!~�K]N��u�� 	]޿Γ�WǗ��ݏ�!~�＆�1L!5�V��
B�1	��`Lu��&ֆ�[�֙W�O��@Al�Q�A!˗�dtٶ��3W�� c��	�w��@V+>2��\�W(�!���t��?x5T(�%o�������ҟӧ�� aZ<�1��3�k*p�<�u��`P(�X��B �Y�Zl����JD0�ّh%��&(��2�e+j(.���F['0������;��Ͷ��rԦ��A�����E	 /�M��}�h��:35Z��Fp�b���;�x䐲�YW�)�k&��K���D�+k� 9{�?gsչ7M�O,�'�=\�i�H�}ɡ"�Z8}�@�:�p��2CpN�&q��Wt�Mwp�������&MN�B�a���\k���n6��5�~|�(v�����O�����ň۽�3E�	6�j�7���C�Y/>[6(�C�"���9�k���\�>#�$�د>���SC�"�P��w�Ș��й��P��J��<�|���z��a��s�`�S��Ģ�dZ�S�7�~�D*R~�����g�*K�D�[%<��':���ո׸qR?Y��/���U��*��pu�T�}��`�����t��<�r����G�x�l�yE��-���"�V�W��#W�g]Ĕ�͹�F�UT$������t�p�@nk�H���F���Ji�(�����6������o�!��_���� ��8Y��Ú��N��
>?��rrU��:՞"gưRW�2v���ߟ��N8��J(�<��4jPOj����htW���n���� ����D���d{�k���J}�&��CF���;�yvu�\��s^��,k�����<� �7u�ev�h��Rx��k��)�g��ɠ�v0(�bSZGS�(�����dd�x���H�bE�#�=(0T`;B��_�u�E��BP��E�dȪ����KR\���#��y$Nm<�^/੅�^xF7g���p 7�I���y�4҄�'&���5��
]o�b�5p�=�R�Ì|N+������ j��0{_<��ί�"�|o�`��O��O�7�t<PM:҉���=���0��*�P����f�����AV��5Q�fV<$��2��=�B�;�C���yЗ[�;%O�g��^=�N~�L{�a��v4l[% {�AS�"��@��mw!��C�C��.�9J�#]�G��F���!�}��"�;d���UD~6־]uӴ�1L��{�o�d�)�,oc�5���R��cn��XP�|���9򃵆a�]�n|��k��UQ(j�g���g�W�XY�c�r��D�1�����Y�+���6t�]����Q�N������=������A{޹���<���,���fT��2� R0S�U�KR��'�0F-e�-q�1����ȴ��&e�l!��~���$��{���P�(�>��3�@ʍx@���I�'1��@K9�}Nz�����d��8>��+��x��R�G�F}AGL/k}4��h�9 ���"�lt�>~�$u���hM�F�͟�B�I��>�{��8�L�p������R��FK3���Ԣ@(N�k���Mi�IXe&�ԣ�����f���紈rU޿X�=қ.�"�8h�V:���c�D����!y[|��J(;SK��U�������7�p��v���b�w)�9MKW����#�J���y��+���Z��S�T$9��+d?J�^6��`���'<N;���C���L��w+��wR�����̙�)�MfҼ�q���Z����� �� ��L,��e|Ti�.	5
�ƺ�	l'h���6���D�r`�;!��:�E��hܼ�n�Kq�|�y��@����5pڤE9~�7mxN��=t4���B� ]�G`w���mD{zV�~Pg'�E��r�k��u�j��u���XR�#!@SF23�K������� ����0�@8�4�Kkv�&���у�Z�>�,��J�Y�0w	IY�V#7�)s�yiwO�h�8Ǹy��G5+�E��wI4=�E�,���s�B��8*t�I7��T滦�oǳgF`QL]n����<�x����':��@�=�JIΜ ;�e��HM˩V�).,���o-�[���5�u�#'AG@�F��W�H@��ě6m�#��ǰ�T�+ew|�x1$70yu�U?�$W�
�'Js]�$~7�Kn�sˣ��хRSN]��z�G��ˆ�m���P�H���!#`25n+������)k�.��7����ͼj��I!��;d+K��,�q���Np�E��m�(���$�l����*qɮ!H��Q l>�-�F����p��O�I������R�)V����Y$*jbqj��^	�ug�5"ė!�ݮ#�E�p��E�:&��,��}���W���L����π��ӑ�&4��Ξ���_���!�Ȃ�6m ք�գJ}{�n�
�����cR�8G:V�k�>����Qh�vFܒD��P//@�Q��
�&���K2�}���q��?dI�^���]SV�>Q)��S߻1З���B�7nx�>M�^�;g8;��g�Y3
2֊fQ�U�ޘ����9�� ���Q�6�ALI9bo���&	�}�H:�w�0J*T3��d��v�F#}�ʷ7A����Ӂ��$��˱�Db�4Xna���b�3���6J��n`�:��jtn_�����hc���d�D��'s�l��B�_����h�������@o3�ٖ��*z���l�9�����L�*u\%�N�u�2,S��~�<t�����q$�tƗ��:�%M̈́B�[?g5�Μȵ�1�R�'Ʌ\�Vc��1���3_��^�	B��h��Ţr�){6/��F���b�'2	k@Sf�4���j=I9Y��E������ǸO�#�OC@I����MJ�8|�Nw]��\,��e�%Q�L݋P��s��2��.�2��@��cl��,J���p�p �����������1��$�wWAaʨ�#{�z��ڱb�6˟�µ�p��Mk˽C�n��Ԯ|��WQ�ElOy�|t#��i#3ܷ�8�K���)�=�`�5�<�I%�#�_�hD^S;5+�z��  a��R��f�t���put��u�� ��[x��缮F�@����u�lr4��+������&��]���;m/.tt��5������m� Z5�! ���4�F�m?h�\�+<&g+l��߼�"sW|��%�?B���]Uj�7	)N3rB�5�s�+�6}�[���INAypd
i]��@��5;����7�Fצ1� �qHץ ��4j	�����d:nFC��(��]�f�?�~@�u�Bo���)�O2o��c�<��`=H7K�oM^~��ly�僒fTK[�MK���.3� Z"��%�5Ҧ�8k
ҹ?�1]�;�aA�XU y=J"��m`b��F"���<8���.n��="�O�{�y��N�Qw���(����%Қ��as������ׄ԰Y��o���iYU����6�9]2��\`݆J�*ci�u��m��6������4��\!� ۽��K{1le�/�tC���\7�2�>x��R����0�%��?�2
��fU��d5���o�L��`��#��@���Q!k�F�ki�^d��M!�\<r��*hܪ=:���?�X�����6"��+s��'��\�
��ى�u�N*��7��o�q]��*��_�� ����2��͈�ļ����<oԴ��w+�2&/6��"�8L�����J<kꭂ�u�����HxT��a�0�L�k(l���cj,Т
��CzRVDD�c� �aC:vY������t�E�S�8���ِV3��',_
��0FS��,7`W�+�� �|.���QE���`����NcY�s_�xh��?+Ͳ�CO O#��1��y���a�#���o�z4�^I��X�#�$�@3��1��i{F��_��Kk�������&�S A\�Ƹk7]��ƕ�o-��ӣ��2������~�9��Ԓ)O�{�$��3Z�>�"}�z �5���SJ�X?t$�lGf�C�����w#p+.g�	������*[�S�1B(+@C
Y� �������rCʡ���.n��܁�.o>/HP�>B2��\H��i�B"L�9W��wK�U��ͦ��Ϳ9Q;c?��g��NK� �_�g�,|r6Io�ij��"�,���*���3�xC�sܗ��T+�1�����b)����H��y�%}�(�}�xC*]���dQ�o�Dn��d��G1u\,��-���)cR��� �J�rQ��V���5+wy�~X���3<B�d!��{�7;�aY �_1-5�7�B��8]���u
j�|�]~�jSN��-������f�A=
T���紜$isk<�-o��J���T�:���\-��H�Tpi�Z�\0���թ
��������u��#YD}���ޚ�+S�?7���Z������&��DR�ˆ�g:h0[���:���D<���<k�{� 0nP��c�Ev���6�+���ȤT�یF$��Q&���O]o��z%F��b�d��\�WZ���Qum��.}g����k�h#��s�U��ga���v���Zপ1����X���4=�7|Ř���ʯ'� �;͘=fhwݪ�D��Px����,���\l�U�X��J��>��XN���y�	ʨ�Q7M�PL��nq&��̝��E����rˉJ}�.k;����!�Dt7"���(R�c�L�$߈"��i��{efyG��h]&�u�D���98?����B�w;]l�g�����Iz��[�h9�]��1����o����G#��6�4g#Dݯ��M�׻L߅�u�I���a�
Z-��P�1�qۿ��H��5͠)������D��'������_�9�)���-]�xn�� �����@�`��h�~�>V��q�hf'%�]} ;ė?�e#P�R�����=u��RL-��Ì��W�����]8�K�'��� �4��^3�®C`/�t��X��Fu��bl����[c�{3��>o��@!�c�B�8�ow�n�6�R�x&�	���[�@-4��U����9���vg�Ҥ�r񘠖�I���-�Ա]�K�Q���ou�-`��(�/�>�����m9)�4#�>��*�)W�D*q+�/+���Fj����� ǔK�Y����a��^�v������]y����l����t:�0K���?����b�h@�$���J�ݟLڎ���R�`��:G2goݒ�z��=�:��� e�t�%BUׅ�H�SÞTH�jb%E@L�P�8����{#�g
���9\1�B�/��k����=kH/�
�gW�q�`�E��GA��'��O�J�è��o�~����N[�[���X�.	y��7W��L ���t��ez�F�s�^� �}Ҏ��P*v���v�:S��Gǀ�g����ׁRZD�Y$�'E�T������9���6(o�#���g���l��ڛ�'���}�m}u�
(����S�l.G�K"���n`��j��:ǅV��{���xޝ��Z��eq��@wq�
�Q$��{c` s������R�!�=m)��6�A�D�U�Ԭ$ ��>,9�-A^�ߚ�抆��V1�����Śa�e����zJ � ����H��;�DN���(ܹ�C�- v8��+b�|Q��7��-z@:=2���`-�ǝK�^������D�9��f������fO6�V�Q�qFyn?,��hI{������ۼ�mp?M$��'�2��;K�4#�v*H�>�=����/��l��Jrb�p�2��"��ʠ<Um����Y&ZVu�k�_�����$Dk���Z���(at��."��a�X�T���=`�<���$�)���䔠r\�����Í$�EX�5���s��S?ِ�+�D�H���2*��E��)kp3=ryE/o�[/��&��'�混��� �4�"_?Yf���������#	�K�����&מ�;�#�Z�,]{�`6ij���e����<�&����a��	��,�?�%����W8�h���q�����!��w
ɪ^TTޓb h,3sn���N���=-�j .<���S0�r��9�5�������1���j5� �Pu��ז)f����`�W.>ȓ��t'��P��� eȯOފ�r�W7O�"z���-�����6*l��
���%�[M'�}�/�q1[6��c�U�Jv*I�;�����<<-�c%�@%��Z��;��Y_���F�>��W����G���<Y�N�m/"I~�f���z�Y/��H~OQH��4X���p�E_�"�#X\�d�l �;&hiD4+u�Ur��D��/�ނ�q{������`)�6UV�}��8�{Me��J�')�%�i�Y����;?�X#M"Җҥ\���1;29�b��I�ݧG� �VH-���_S�{ a�r}�C�%"�dw���OBp��6��q�xg�`GS���ۍ��@|�q��>[���[&���v���H
��[��7~�z&+e�S16���F���»��Oì�J�F�"��\��v�ʒ>�V��8PO3�cQPLն"Z�:��1���_�$�-����/V�k�[�b���6	fu�	g��Ԋ�o�]����Kť�j)��H���Ϻtk���+�p�m���v��Q,�s�{��hVo#�y �LHa�f��%`"W�!$���W9JWHH�K6��% �t#{��3�xؠP�5��8�q��Vy�t} @ D�n��ٟ���"*5;s�Q�6�,e�	��ceԲ-�P����� B�_	��X����o����{�z"���\�."S�\�7�)d��<��+5j	��^un���o�G��lr�wK�Z���c�$>��wb	R����)p���M�(�k*7tT��u�.���#�!4RO��	��R�L��U{'n����Z�ŵ��0��r<�W?�Xs�f�z��`����j��*V}I���.��)���}Թ b+ �Bt���%����Л՗F��3zD�f_ y"zZ�p�X� pS�����A�,sͥ�����Yf6�?�M6���-�O���ָ&y�),�$�0J�l���6Ϩ�6�����W=<h��H�I!Xf)҉�.1�c��i�URd���
|�xJ8�Ǫh�rI��+�]��3�{�;x�u�0���0��ڼ������w=,r����f����&B�&-�ל$}�3��/���R�HM�D@ݺ�+Wu޲����w����*P��?j�엳	�:��g�A��U=O�j���C���x�
�wA�p��m��r���u�r)�OcS�(@��B�4�wJ�[�iTC/!8�̐�q��9��bP*t�$:Cr����^�t�Y ���^.�]��s���ۧ߆���7$"k`����M��L�r��JC,W�f������	d����F���-h�̅�L�a��(�d0�2S��?8�Ӌ�ad������_�K�� ����-5m�S�eϐ��`�'9'Y�\�{^���5� ;EsΰD%h��&���"]���V�XC���a�TUL9�f��~Њ�W_T��32V1��I&�p���[w{��Ƈ�bga�+�Nrg����"z#��;��-=J��)�۵I0��̲��	&֞�v���|.3�|Y��NR�6T��闍h'(9H� ���ŵ�rKsӌ|���w[��W�L.�}%�fS�=�~��J��sS�؈S���!�50*K��sR���W`�Q+	��u]s�
��Y{���Nѝ�f��4۱�?�����p���Z%��?X2��Ŀ�.�|��j"���ц�v��xD�K����.O��p���M]Լ?Z%�(�&X ����:>�~�;oL�����co�o�y�,��c����U!Tv�h�rj�6�Dl_���*�zޝ=��M;z��G'K�p�� 5Y!�@J����H��:��
3��1\��BH0�І0�MV�X��Ӳ�1]"|�U
F��R����	������pV��0.��*����"ש���ݩ��#F�("Ŭ��1ȡ0�ip��Y�����ːbƋ�b>;��V��ݴLw�0o�@1٥Ib�L�+wE�E�v�ŌH�
��+���m�/I���B$��	KĈ�w���l�2M�#֗�!O�#y�ggL���R��x�'I�����:?��'��xpeA�-"g��� �7a`�"���l�Y�O��x��C�eHo!����&�}A5U��۱�#
oe���i��+56���L_�����i�gmUЫ�N�e�����Ǒd_�(=F��:��#��ge'�� >p��Y�n� �3����T>��X���Y��H�E#�Bo����L
¹,��\{;~�le5
�jDL�>�\R�8���#�'-w����u�������ة[E��k�*��a������ED�Vz	��
����m�ۤW͝�^ޟ+���.[��-�RV�畹��^��^�l��d�Ik��:_���0��ϭ����%gf��GՒ�ç]uo�$��@�v�9�D:{�n��g�����������,R@︨�+�紥G@1|[c�hF��}l7tԶ���q��$��PN��� �#�.ڶ�{��S���z#EpeC9��ڈx5��c~ y��!��m��o`�w_�����R�bhJ��5��i�ePT��Kh��9[2.�Z�G���2F�b���cv�؟1K�Q��.�o���j#j�b��uƕQ����'��Gx�8@r�&Lepz�7ظ������%6���K�)�S��ɰ����Xu��dk�"ѵ<�C#����e��~����m��ֽ����je��F���X�ވ@�eN���e��ǚ������A�`G�I�6(6�ȥqbl~t�Q��Y�ހ2�k�t5�K(�Zx��3�J}�Q����i�����0S)*+�њ��$��ӳD2��O3d����9��#�x�8�P匃��K��q]LhK�S^���I��z5@������<n!kT>;����~���yoG�^͇����h�%���|.��0�m�.N�ʡ_�y�4D�]_T1� �׻�[��}K���4y��v�җ���C��ES^W�H6����4��'���*�q.��ȴ;
Y�K ��G�MS2���ƎڧdD��m�t^���{;H�"N��&k2z2�r>�:�x�u	��Uyw�0W���5g�:C�Jg�e�{fI���=V��C�.n��~��J��>HI�Y��s�~��!=�(kb�����GH����Y�W�(S�'P�AE�:�i�?|�Y��ct>f �@�6�P75\6��$z�!misj	�e�I'C��@���`e��ӥ%@,��`����P,3N�[��v��(}��s��Z��J�V}1ڰ|@	��[YCCX1�bq��wq��X9�"��WNA��ʇ�c6~�}��0�r�|��^��z� 2�װ.��=Pu���7�#�	�T��:��K�.z��.��o�[����_:�	�zt�Y/D����]��1[��$�J�1,��Q.���Tx�ս�%!����4WC=[UwB���1t�}�fA�|?�������uK�O�8���;i�vObT�����Bf�e h!�����)n���� �ڻ6�+�@B���\��	.��9�K�FH+�TS ����7H;O�c���x�R߁����������a�<B\py4.��K!�L��z����^;��ЊU���)���7?��V�r��ޮa��`5-:�_g�J%�0�)'"x2R�Z�W>���( �:�V�i�t���4[�V��+��1v(��y�A�7��D�I�:GC��q�a!!��`{��z������J{L��9�y�!�zVy
�7�qǚ!\
�z�������o�ro-[�a�9��8��Lo�
7Xp<�ɉo�@2�5�n��/���;3f�b����v%ᑜţM�0ҽ}�� V�_|��0�q���d�:��kِK�2�+K�����̎������)���������o8C�u�������ٙ6����w�����S��]�xQ��p����Vt�T�Q����YI9x�T�ke@kZچ�љ�S��脸��za��z��)JP�b��m�� a�z4c�/��[U׾C��s��	���Κ+~\�as�	�����>��s�MA從?P�zOjR9;�8>�D��|�^��o�0x� '�8�DԂ�ʵ#��f�o�w安2d�)~���#��Ð*�凞�iq�8^�|C9cЕy�����PR�l���q��²��@�D�W9�t�S�<�L�Ne�ad0��� 0�̫���J���>�hA�ѝF�U�Lh��sؓ'M�zς:���'��8�4/>�J�H2�Y���@鵴(;���W�&�)Y��=�@���K�0]�,VU���_$Ӌv(�?W)?�C�x6se���M}����`�v������q�w�¹p�9�h]��ԗ�vcMF��S�5Z�r�b}�yh�ɯ�C����\�>���*����孔��V����#�� ����jiR���290_1N��̥�⚕�3sUn<�s�KP$���O��:C�}�JT�������*ۻ��M:�fߓGa�qe�H�p����t�i&����ej�:�1��y��k}rNDދ蹴�L��92>���+���*K7Y\�i�%�J��Bq�~g ���1V�|�J��;1���Jr�❸s�"�;�1����,g���̇I)f�<�F��pA;��fM��B�Ÿ�J���D'J�G�:FM!�P2bssN�A��.U������ڕ����`L�.s>�=��T7��^@�LQi��
�ec�S���������r�ʖ{� ���� ���Oo�+�y=��fHlVY��IZ��2u�F��ٸ�M�Qw[=�/l�}_����%��Cѕү�n�07�����qp����u�~X��#�6���m�`���H��� 9��9
�����2�p�W.�����"�1�{6�k��f���!����Ai��F7�F�D>�b�q@@X_b�C�O���������N���=[5�oQ%ʸ2��zq���N���7l��x��.�t���>�рR!O�|���]��pKa@�u՝�Qb��Gt=�gHM�$�Cp?UgCkK��E�~���_V��mnJ)Z����-�]$�~ [�@�;9�Wڡ���H-�b�ls��l%�F��?V�Q��G}n�%Z���v�f�"OGd�n��B��x)XJ4���.Mu��C��gu0�m�Q����|�U�Y�֧�a$�}����r��W`s��ÜF8q�+)�۱���=�g�Ws�[OS���,����i����W	���ܕy7��C�`�o�n/bT���<M�>
?�~���P�Č���e&���P�ř�9��O<�g��W���X�v:).'�_ e���kr��h��]�`��g)�G�l����9��)���'���(_�x=�Nd��F[<x;0���eh1ɫe��z��Z�Ʌ�+���O��V��qRum�:T�q6A�A�����9��ag���e,�dҴu��DZ�S���q[�����)Ų��� �%�j�aKtQ�'�Q�b@�Ѕ�E"��lg��q��na8��\�OS���#p3�p����	4���܁�Va����}Zv�*7+�	�/� XT��G��Hi>"��Y썹����\��������6t�*����?'���<`��.G�i�d��J��9�i-��刂~d�����v�����P�=�i駜���ҟ�)�\Wp�}j�UK6r$�f|�<�!�2����>#
(��a�ߋˢ1�<[�
a���|,�Q�����7�a�G�ܐQ���f?�z�ZG�|s]�4����'�:��T<;Ҭ���ɺ�M����-�J:8V�nkj?O[�^|��T4"����F���}�:��;�����	���g�����ݮ�c�3Da�+x�&��,su�=����b��,�E��_Xp�����b�(+��]0�M=C������k�Lqy�4/�AA"�캍DD����~U!w.�\S�E?�#��q��R��\��bDOP$�De7���]T�9���=���y[��ߝ��-@�*� �C5?Uz����)�;fdx�vwlJN%
ә����Q�ޘSˆ�M�/nc0w�&�g�a�1�t�+m�vN;����(�[��Ҿ!g���W�����L&��0���I�Hy+	7��+Dm�j{�ןk���M��!7�~t��:*�/�#���{��,U�-&D��Q�T�¶-Bv+�l�����o����i������;��ʁ��O8*j;�� K4�Oe�'`H:A��
)�ㅘ�懐��dYZ��u[VU�9|�J#O�Ѐ�uT]0�l���˃*��o��c���r��<r����%Y�},�,3����
���{��.6C�M�ՊOV�����Z�7�`4�MuPY^\g;�F��Q"��w�2���#��5�Z�3ީ�+��m�"C&�@x+b�}`��Ĵ�Y��P�~��1YY:�L�������X��&Z6�櫣xɀ��މ�c|�M�Y9'��|`C+��e�H{�KB�O�@Ff��Ꮆ'���#'J�A�����Ƣ��6	�+B8h�B��R��� $p��&n�
��iۃ{6͕����뤵�Ӹگ[/+l��]�-���o�c�~v��v+lx ̃k�1���;N�2��^�
�)�黾��r���5/��d�J�B���U���+��l+Ҏ���aJ�f�4���[B�6�]�CT�����m���u<�����;�ƈX���M��h�S۴�fn�U��_*�0k?w��>Y�Ma����6�˸%�Q�������nS�^]9J�`�Ȼ�6/�ܧ5�$f�\T���ן+�������,�F�C�>{�OQ���BwG�sf���}p%ѫ�$�+�)<Z��`K�Iב@?,�YF�<��CPMk�<��,!T:I�j�n��$� ��وQ��Qw��1;Oܩ5�����H��O�qIs�� ��r��W�S�nX6��]/M��n?��(5
4�3ĽRn����u� �@b�66�Y��p+����uip,8n����rT '�0wx9�~Kߜ��4���0���V�`�UX�����	D��;��ܢ'p���LU�Rf�wp҄��~�-4���������JQվ����[B��V��w���
�ALn�mmD�����;���u�A�兂�i|GKq�o;Q48�T�+�}b�c�{�!��f���X�:����L�������o�9��\a�K��ݰg���EMҢ��L���j(�t�&�oZ�+j�pj飁%=]��gF����04b��-�)	�����EW�7W�F4�d�}���j��[�wz�_H���2�/+˘n�E�`B�U}����8~�S����&¤V
�x�Q.�b\%^C�H ������>C�f��w<1�H���_k�v~�H��m�i�n�6}'ű���K��׈��ԗ��=�$���|R��z]41�$?����0�8�O���P�}���K.������o����8 w�^��4J1|R�7՝ލ|Y ]�	��3��x�����m^ȓ���)�*��&�;�?�Z[���b���H���;�Mx6�r��=F*���2'����*��C�h��Np�o��p�'@Fgj�9&����z�&P(7H:FM�?�:=������c��v��*��؊T��1�.21$�;1�0�����u��E�q�˺�͗P�[��:Y��(V��{2V!F<xL�3@�C�9I�!%(l$�OM"4�<�S���ݑAȞ���1H%��u�a�r�� ����4T����&!��7�X.A�E���'Mr�ը��F������� �1�Qm~�M�p#�J0?|��dw���ʢI7�M�u��۩���B���;Gd�f�UF��儛P�6���m�����!"z��hF�Tf���1��x	�&A��g�K"��S�����n�)>��� a=���h�B ��@��	�ye�p��;+���ą$3�����k�z����W����&�|!���q��m���~� �uf':�e��G�iL>��c{l�&;u�ܠK�@jX�BE�,�zGK˽��%ȏ�՗P>l�-���kQa���f��=׃襽��?� ʠ����X(UR�mu\2�<>,X������A�3i� �F�}�vf+��e��t���CzHZZ sjq�������^(	�����|0�%�)��g�/%\�Rl�+����˽�bD.��r���� |fj"����|e�Fr���-�(,\�#�w�o{ ��S����ºy�z{��Lgg{��t8J_8��H/aGaX�S��r�R���Lވ�[���$�H=���'��rD��1EC�˫2�����#d 'Bȑeooެ3�ia�<�)������$��L��%��q��]O��!��~�� �&�����Qc��q�U*�����tHt����H��#���5|РHPTt���������+v+�6�����o{#���,��_ŗ�v�η<W�-4�j��ϿF�,YouC�w�:'�o3�Y٥���e�8�5Jpˎ��~�7Kӂ�$i�����<鮤�΃��7ԡ��{�`��Æ�Hyl�ĹH�����w�١�+��M���"z%$�)�m[d}���=�u�|�@����6� &��B�!A�j88��y^M���w@3��y�:���}e˙��ҍ��pXH>�r[��%����F�N��c[�Y`���������l�6'=������XO:]Ē�<Q-m��p��F��b�kx�����q��97%A5�!@��� ���-?�[��%��FU.�j��I���EС� a)�����5�x�=��T�Y��!��	n����!^��K�Y��i���#�	����(͛	9������Rf|�m3�06�W0�V\�'�5X|�P;�� �Ůj^����3>�Y�4�T�����e�H�dC�i�Myـ���\���Z�1i��|ʄZ�/KUg�JkKCԁSE	��䙨��հY���#EIw8�����cQx4�&��B�Q�g%�F0��ÈE�pi4S V1��5CI�a�N�#�aM������)`��Q�`󳵥�r�#Qz�/�¡����7�t�Q��ρ$�bj�q�ˈb�2�YO���t�_�}�5���S���ݥ��8!�h>`4�Mb�˝��~8�>�8%�^�[� ��%m9d�0a��![h��'�͎9Z�v�彝H����d�fo���cnIEK�H&%�֬����4�@�'��n���m�����Ж�ӗ�X�̴*����u=��t��0�GM'�|L��,{�|�����oq�q�S�������0�����J��ya�[�&�֫Hqପ�-�,�㱄�^�+����([7m���Db��۷��L�'�p�0?Ϯ��m�|A��/,+�%d�,WQ-
`�6~zG��덧�s{�݌�:��~L�TP�+>�5-�¬����� 'G�+}��A�zR�{[�*6E�r��wݗ,0��y@�	b�r��Z.5�jl��EQ�PC��:@�<��e�<��`���g�F��9�mn�	A��ü�hY�z�$���уɁ%~��n�?iJ5��$W��AԊ�c�G�T<X�5�6����5��A|� I��	�U�;MS�&�N
���s�W��x|,q�����A�F��f�4����c4Y���E�5H
vpPw��J�_�$1��ė�@�=��v���R��X10�($0��vNkf�&ZYv�im�1]G�}oZ��ܧ�Xe��l��M�$�K(b�Į^Vqื���D�$�kJ���<���O�Hn� %9��Gװ �c�.��b�<�~��_l�귂GW�&Z�/t��Iʪ�M��Rt[�����R;-?qnx4�5OP�����xa�.dㆍ{c��s�� �ù�ўޙ7�����;<�H%�}���>�V!��������J�qX�m��c�q��RvD�:>�<ͪ0��˥����ɫ��@�a3�@����O7� }ʏ����1Q�=iZ
t��"T��JO���%g#�Uj��ߘ��x۞�]��=�"��/�UX�^�U�e<��K��|��w�N|�/^+�-�Z%���PJ�	_���+���ǻ���H�M���]Ӗߣf)�����T��̿di剭�5X�4���5��Y��pI	��q�Q��l��E�e��F��T�=wD_¸�X�tH�J㐨�d���ԘT����&�5���F=�Iud�rP�ؖ>љ�訵x+�s��lӗ��Q��(�(���s���t��*6�u�f�J/�����'���j,���1~L_J};�}��V����'Ք��u�j���c�Y �y�۰G���H�۱&V7,���9��W��8=�/S�z��l\��o1�)��I�e�@yv/o��9�,["�c
�s�7����&�HK��z��Bsh�~�chD����~�rT�N���H�p���$�Љ�ZSi�������<w����59E��`8&�=!̸�}^�P�EJ��7�s�A��{����uV�~k	�~�B�@!��}�0;�F���聩��&n�i�����C;<�	�d4�Z����4�������^"ɟ�+�=S�9ƴ �Cqnv�	��V<���a��v>�Z9V��^�^ 1�H��,�����E�qvUG@l򵱟�v�@�	j�����Nk~��\�?<l��x��"xW��Oȇ��Yrȯ���q;&��������<�Pa�;�IH��IE3�]��j�� �5F��\|�lz����([sK+�D"���B�8�g����Sa$n�c�;%��ȢF����^(�0r�ҒZp��K@Zjg���yI�XдP��fj[��������A��ōa�Cպ'jR�B�ҿn�Cdrؠ�=_��*^Ϟ������7mN�36�i��S��K��!���*d�����	p�����π�;Q2���	A
�	��h�w
�Ҏ9H�`D+R��
�Xq���r?��v��{ђB�f��ȦK�K�X�A~�
Gw�ۗY��	������W,۹sɽ,�Ϩ�?\*7�?�َ�{��}�+�݁~�):p�XXx:tМ�`٣�4��\��٦�G�"��A`~��y�P:�q�$��"?�<d3�=�iG�o7a��j'ʺ�M��8	�Z�՞ b4�+'���
f<u�2��D���B�rŰ:[���	��Tp�n��~2Y��ÌA��t
���f���[��v�~�n$ž��>g�������dV��z�x ��`���(q	��X��~�j�w����z��%Ӆ�O9�I�fR��8��f0����]G@����=�#v�eY��dA_S*@��%+�}-���Y��� �Ҷw�gz�_��������]���9[^7�n��jX0��(��3�����iV�#ӑ.����z��:#���vQ�!�R�v�s�G�k����wPݔj*�"/��kU4�b4�皷_ (����R��0�c�Pt��D[��m
�!�x�!���|��C��=��V���n{�O��mOrJ���q�3��d�!7u�����2�+���3<��O ���*�4.b���v��7I&_S_A�5�0c��	��_��s���;3*�w��q�YW��TKe(|�M
�'/��'�C�鱾�AK4j��N-�R#�����<\������3�N�a�X΍<�z0&]��v�^�Y��[a���\7�[���.�͐T� W��p>��lGN-ڨJ`��ar��p38���M��C�Ѱ8h�"	�)�\#2�n��DP�/���.�)��j�W�gR�K�|��;ʆ�!d�����9F`�Z�����w�5x�ךh�ۂ�zMy4��g[L���;���؂��i��W
=��Œ�i�\�I鹁EW�
�d��C�p�oST~�k��@�a!k��F8�~��;PCLv\u33	g���U�D�i]��v���5N5�Iɸ�8�"*l���z'皗����'�R�I�V��q���v͆8���Ixb>�N�ӑ�먏%0�N�{��@���?\ݣrJ�����PK3��E�NE�*���	bz8'��NlN��S���E:Ҋ9/��(^Q�]wE�	�Q��U�R=IU���Y�ܲ���D���h���v����z��U"�o{�{�������/��M~�<E�a�y�s�{��K�Lw`�μI��r(�G�[�1��>�� ~�1��U%�U�}��-���Qʶvwy#/
�R��1�K�����z)�ۉ�%��6o���@{3˦��"�����9)K�.�=9U��VC�+Q{��l+����x�ނ��(^4/f�`�)&  ��o��;���v�dC�Sk�nB��1�d��^�Q��ǯ�H�17���[a���Y�,tli��G['g^��Ї������UC�
�f����x�	T_E8[ �y9m�c�QK�����-+�-�cf�ϒ����p��XƐ� �����g�]�A��
��1hƏ�a>��<�v��8���u�5��6G'QT��g �k4+Y�M G7��� �͎w���0���Z$f����8IH�>D�Z%��7�G2&�:`lњ��&)��Vɂ�^�4g��g��Y��3
ީu��ǹZ��;�'���DYDR�#ՠc���e��Co���&��EzƈVd�Sꗊ��`� �-c�"�n9٥����(�Ɏ�@��J���F�$�ۓo�L�~1߂��$c��Q�_VE�ɧ(��Uci�/�zs�HI$���L�?0��0�����A�V��9����vCQ��dM�S�'f��-�����?\	������f��G�j���q)���m��5 ����r֌vA��ӳě3s������iӷg��K^�|:$�ɝv�����#qk�;��qCR�v��W9a����e}��1�U�Ґ�w�d���qȲe�u���mfJY5�&W���P{1
��μ���n�(iXIf�k� M�S�sxJ��;�!vGD��1/Y��ZJ_Օ����"�u}�ǡ�&��	���@�,��}ir��Z��&�����]S���`z���u
���`��wC�m�8�bt]M���W��:������eW�;S�Sݍ.��"1f��
��v%K�=h�R�F�敘W�eui?_x̳^|7��Upx��X�\m[���=���]�P[Q�������,�_@�ۆ�;c �� �P 5�;��q��{� ����iɉ(�#SA��.����3�[�V����a�be8�T�/5�ގ��j�K	�Gh�6�[dH��'�bm>P��Q��J�KUB)�}�i�����bl:6��C���{��H8ұ��hr`�Z�-#aY�������:���'��`P�_b+���6ϰ<t+�r6pw��ڿ�n�!i*_��k-�K�6)�D�e��ή��~��!F�/ �U�[�����N����}��h\�n5�*H�GC^9�G/(�5�.,1�Y O��^�#�`,�+����G93a���P@9�ƕ[�|��k��I�)Mq\��4�S�⾮�����A��2�Yw��X�8���Ɛ���a����VG|x��C~��zw1-�[�]A�����E	0���/�ұ�6����w@>y��H|�H�5���}!�{̗� k�SY��5۱�A+uud�)��\[��� (&��猑�X/���B�G@�J��	���[�������·M�N�04�G�8%ӥ?3K����㰖��e��]���bFvZ��+�� �*.[��@�$��l��k�i?��c����� ������W"��J1�ַ۔�b�}*�Cʁ�	B���G���i���6���U�a��})h�M�I���O����ǀJ�����j���jqB��s1��#*U9%Gq�rޤ����I���u���RXjL���ˮ���P���)���y�A�Kӡ�֞�qkhx�(�`)F�=�#2���{_{�gJU�)��
x�H��ǫBJ��d�j<y]R��'wh,kG�g��4�/A���%)I8y�DP�\�Aa��!�V*V�c��xX[��\SfbJ�>m���~L�������X?�9��y�d��e�~��^��I�*x���5����.���e���#%S�����`Ӄ7��>����������h��`�/a?%6�9Kkf�x2�M�a..�겶O�J5rI	T���c:Z�����g�������BRUI|�R����L���*b~�M�\�:~��0ҝM	%����T�C��U��x����Ĕ'���PUW�л��34�[YOr��'x�1(��Lmt>��9��{��{����a.a�lͼpb�5�lH���Dn�3��5厾�MU��mr8@Y�� yf�̦1C�.��"38�5�`&;<��b��y��)
˵��m\��d�uMG+7Qy�by������U�����஬k�|_ը�]����bG��$5��߭�-�o���93��?�ù^=}T RٝqЦ��}Gm���eEn�����-���v5{d�b��~[Tq��_���E�3��?R-����eC�'����q BJa+�7�Z(�	��� ҳ܅C&s�6��1����&2����q��+B��iq�8RpZ�
vޗԂ��c�r!�� ��cD���ߚv��m���ޥ�k�xPڝ�3�S�8���+V@�4�c.��#�l��o\)����Z�܍�s?(Ri�)A8B�o������B�KJ+���"û��TX%��CeM�%<l��-P�����GT8�[h�(i�_��1�M��~"[m�Z����/*�EQ�b���eo��	ϖ_D�P d���w�p?Z�P�����7e1䂀=�p�4�v��*��V�Ӥ(4@ڈ�\÷eRd� L�-pQ�-.����|'ٳ5������$���/'#\���-��d���N$�����^�jD5����X"�e�@��л�P��e�_J�M��^�mEI!��)^%��S�*�V3ng���ox,$}���f=�yӨ��b|�K$9�S����3zF��/�Œ�"�8J��D������f4�O�SÏ\�����;��D�����O���Z�Y&���<�2ɭ�g��2[��jY������ �RL)C��#�ւ�؂(�Kw-m�Ψ��г��J0h�9bY=d��x�t�V`}�m �o}ֽ�%n�_�'���%Κ��#3�L�ѫ�K��\9�������BY��GJTᐵ{�T�����V��	fv�GM�	�}��M�҇s~:Lv�Cۃp�[��s�{����+q�@2��Eno,R6�����c��g���8���o�$��6M�v���1�<�S�7@:dW1c���G��7W��`&�><��U�5�[|l��g�i�ZB�T3�(�.��B��0���^���� ��,ƙ�.�B/Y�{�|E�o�n�"�l�,AOmd��4ԗAv���Ÿi<�2����E��S)��Wb�q#��mN�l�"NO��f��f�aDo(���I�8w��uj�� ��Hn$a��e��[�V��۽��(u��:p���~���m��pN�o6��J}=c���[��/�/��kN5g;	�`�f��h���w�����rFq	��q�o��B�v?ѻݳ��7�@���,�`�H���1�E��I��krA$3���!	��D��?ͽ{T3=}\���(��%&8���L��_�$�:�"F�)�*�x�×�/���8��nndAQ�������r���  }�N�	Kò��KL��\���=a}�Fg��K@э�]�#&$'0����N�� ��-�֡$U+����g.ď��!���R�/]HX:N+b"��ENlP���cfO�D��hS���M�'��o����^���Ì�9��^��E��]n:�`.�Y�+%r<�3ubχ���Z]����)�o�&`�zPY�T�#�!�y����ヌ������HS��󯱢](�i��:��j��<g%�!HGU f"�B�#k&=�]+q(�#^��vP��叄=O��o�B/��W+L��!p��{c���ދ)t��%;�v/}E��������$a�&��L�/�2��Ě�?`���L���j���u�L��Ō����!	�)��	3��z�+S/d��pG0�65�+�8���v+kb�+˟�;0�W��Ѭ�<JI���_����y ����lC���Ro�[!��'s��2����7�p���_�+��ތԔ�� Nhd�����p+!ֿ�� �\��x����*�
��;�Z��z,�|�,	����g�2[���
b��?Һ����}~���M���||%�N���N)S��a��k��#`ݚ�[�����?������Z�ˁ6��3u�Ӣ�YfY.}�d�����q�ݯ2���(f�P �JP�����M�,�#�cu��k^2]6�#R�M`	� }^'���9muGD��p�u���O��Z~�(��QG�A��6�I"���<}x���0�2,XV�ȴ:�+�Kskʅl�����6��,%B��)�(�����y���T0(z�mS���]�`�&j�J�[�F�9^�->���-I0]��`�񃗜-���4i�i��E�zQ5�fd��w�1�7R&B�g���A:¼1Ϡ���_S�n_�"����LFLo�F^J�P���È�%=0��y#2�?��Q�G&s�Fe7���#�&���ֽ�w�ڄ����[p�Kw���ۮ$n��^�C-"	驰w�R���%�����H��(Ui�-�5=Y���7h�#��n����c��6��'I��EA���]0U���;O�#��7��I�r�W���F���֯��ϙ`ѕ6|�p�'1���C���e�순y6��uc ���й�fU27��*�����G���޷��g�����]=�!f�=���_i����:�a��f0L��k���唀,ؑ�ܝ�)n' ����Y�`}�8��oJ�4[��We%v�[/��j����T��#�r~�`�}���G �t5X��F�5�I��F�m��勒u�Y�{���u���W����"���L5���D��=ޜ���+����-'Ռrlm��@|��<�,N��?���͘L#���b���t��>�WN��';?�p�ۘ�~bş��@�����d��0��ؖ�# ���%cN�c�"�P����x���R�f�Ud�R�6\�m�{�S>�>�L4]Ÿuc�_ ��k-��]�x�so��.S��QM`E&,!��j��L�9B����
{s�<l��=�~@�� ଞ.��	"@��c���j�����`Wȍ�-����|5<�9��P�$�b����V��3��<O�d?����� �!�����&��h�
]�X�wǦ�'fx͐����[��HO(���g|q��,G�v"!Em��v3BJ��|��(%ل�Hi��f�6X�{�;tdt��E��)f��,���L��C�ʅAs�J��σ�-�e�����Ѥ9�~�j)�.�/F�S}�]�ė{�la��r�� �M6��D-�D�c������W��J=�!�3./u>�A�	�\A�X`f���bs��Y	���
ģ�����K��H;��E��&6�*���ip,�	�z� ]�MS��a�g���#=�b���U� B�<D��^��$����crS�踧����M�dU"ڦ�k2����r��;a�;�V_� iTd���(Ll�������C����mD�����-Έ�$rV/�w(���ޮ�����u`Æ��|:D�]�[�Y(=�5�"�����4W�!<vB�R=� �Ȍ"�C���̊R�~#��&�2]b��ȡ8��qZ|����~ߗ��Ω�6*�{�]^7e��j��xH����Hԧ����wc��դ0��ʊQ�\!矵�/x=A�fb�����Ɯ��h�k����"Lt}����GGg���t-ndbYQ�}�[�8
!A�� �;0I�w�I��mE�D� ���;��d����es֠U�Zژ��u��tځ��vgל=J�i�6�*��)w�4bhq`��$L`�'w�l2jI���񷦷��7[͗~�qk���0���"q�+,��Ec05���^�\;gpu7�浽�!p����m�E�����?�GRF�r��#���	�l�#�\�7�~'_?!
�UJ�+���GC9A��
5j���à-1 D�f�5/$N���D�٘�z#�j���6~
�<5����{���*��W��N�L�u�6D���t��3�d����r"��K~Yڬ�@/�+h�dS�9P�풾eMkj�tu7�)W�n�a*9��=�M���򬌉;����<�>N[:�Ж�
������F"v�ZO�2��c���5@����g�5�Z=of��5���G!g�Y��k�S�����Gx��P��p���~�"0�[	��{?
ξX�B��7��7�����U��@��G��Ч����*��~e���?5n�25�7�Ү��lg���4#�aq%[�\=r�e���Y����|ʒ�
�U��qw��t��K؛�X���5��K��8yicW4v%A���7w��z��V{t��.0@��nN,���qb��h\���Z��V�EL.P�w{����Y�6sw� �C4�!�a�{{�M�;%��uM@B�����LZqȀ����(Dg��0�C#Vɑ`���%0����ؒ�CcoT���6��on�M�CD��Sޝ�4,#��[5�|)=n�ݜ���M=�2���~5р�*\�]����]��>��4����msȔ�_ �> z�/�p�)���*P��f�x������_;EC�\��"��9ّ����d�k�`<��E�|�[�4-��%�a,@L|6�MI_3��R���6rU�x��9�a��3u��X��n1���J����t�A�)s��>ӰY7y��2������T�O<$Y�V���yr�(C9i�'���E9]YR�;�4�e�6m�]��e)pe��3ۋÓ��[�8%�"a��u���6XҎ�G��9њ-eM���?��&��>V}m����*�j����|@����/�q�+��a}�|x���i�NO�w՛u��.�<�������GL�7Vvj���$$�t�B� ��3�j�d G"Js�A$ɨ�'�k��dˈ�W}w��O�^���sշ�9�>���m��ysjDx�(tRL*�eT�H]6с�o%����暷j����j����0X�����#�G�\�N+H@v�3�7�&f~�"�Z�(RR��p�(��#,N�ͻh�R�<�}���j�p����&1<��q����I�͙���|>�.�]a��?�g��H�����6<^atX�_����b0	������\w{i޶4O�����N�wݰ�����V��*��c�-�R<�x��U�t[ 	�}���Z��2Xj�[�
��h{����jjU���|�&��eú�R�N���?]��d�UȀ���?�����W��� O�6�����a�uP�JqF|a�1�܎�����g���ҍ BF�]�]6k<�:�@���M�%��}xt+��ũ��>���5��ik)G��ò@-���" �L\��c�������gv'�k�8�r@J�$�s{��痡ž�$�b���߬�*�	*���OoLhcY�ي���A2�03�rG�p��~���9�ۍ�M�(��Hz���������#1n#�;���m���t�B<39�@�1���<�=D�^��O3"���^L���\�Zr��������A���f��ˆ&퉕CO��Kj� ����kM{��0=:_Pb��e̘	UD��@���f��9�#��c��o��s#|���m�K����E(C��
�J��^���+L�/�șD6:xN܌A�6<T�|,��>�L��Y>�z��p{��@�����E�����f���d=U�O.w�M��儖�=�$E|!�Ms$�{ƈ0K�5�xV`����_�8�A�d�L�<K��V���]P�m���d�8\��&&ք v��]@�m�$P�VXv
�*-d�ё�vK�k��p�nd�����Jֺ��{����t�?�F���0���qN���a*�Fǥ!����q��O�@�AL'���ڍP^�]?Y(���R�>��εsv��1"�� 9��X��\ �u�-�<�@�i��/;'ux���3l�p�R��&��y|6�Ʋm:ک�|I�����U��S��Icc�B0P���� ��#�uK���q�������d�ER����3C�7��\�W\��a<E�O���ؓ���9��<5z��S	uq|�.iZwt�(���}�"=����f��γXi�VW���|���ρy�,g���5s�Gչ��3^�3|�f��$j��ʩ��6��Κ�/Ʀ�|�T��|��*����I~�%R���TI��+��T�(�Ʃ��Ƴ�5��+����\H��3�)=��Bh���>�~��/��lC���> A�b��yMs(t��wh"�rJ��5tI<�/�h�E�^Һ��Njb�]���M�#�<�Ӌ���{ʊ�hz�����������VwԈ\�+��g�!q_�[��f[ �A��5�Q�MHK�А*��A�u}��q�H��H���:��h���}r�ߝ�q��<�^�c�ꚝ,�[�
�=/���9�v:u}ӱ��;��s�n�d��(2��Vk�u�9i��l+�9L��Ŗ:�J0�Յ�����j%@���׏,Q�3U�-9ͤ���7�,4��@����ʿ��fY痉���Z��&��bc��+g\�^`�&��� �d�/�`����=�zk�,	|.1Ft�r�����sqM�|ڏ�ni�gA��}�A"�.8<9~Af���r�*��{�G�:�r��Ɨh��˅�������#�Q*H�f�'׬1�Z�%����X�X��3*���1��*�KkPI)�#R�� �K��_J��["▨��C3-��B��ay��@��-:�H�7�"^����O(_P��ه��I6}��\܉�ʼ"�����D\�xÑ���͊X�p�,�P��m}�kmw������O `+0���H�h���VH�ݑTQ�	��S^E:I:)]�S����P�
�I�
����� Y/�&0n������隨V���[���?�̹K���h �M=\OJ���f2��Oן/IY��a�� �'�-��p�ý����t�&H�Q���]�(�B�R<�1���[ݭ|��$���,+�E��߿3��O"�#�7��>#��jQ�%�>��6����wx�;t&i3o�Du��P���:TQ�H��]TDB�0�F���4�uD7��?`0�������&�	Y���0�_��Ύ���1Co�Y��"=���lӃ�r[7,U��ǀ��J��b{�� x�u��Zc�/ ^�gT1:ϖ�� Q�^,~�9W�������ӂl.�v��Yk�8<(�Ţw��C��(�E'!��W����j�i{��`��d��]l��u 7��L�h���8����H��u��.E�+zb�$z���JK��L�:�6��2�½�5�|4��e��K���}c`�Pu�ﳁ (���[��{�a�8=�U!���U���y����n~m4F
q��`����\î�t�{.{V	���A}�QT��(��ˁ�j�׼�bQ:Y����FP��h�<�
���_�!�-GԬ#�Y�#C����B�̳��KD���~.�E��L+x�\���$�-w8��AjeR\�}#��T5Y͟3P�uŽԥI.�����
���g=r�YS�x��a�.��Em���~Z�^折���2!��fϡ�� �4�"D�k���O2����)n�xYT`�5����2�U��ݛU+���!���LT�t����;:��Ftx.~�����$�N��<�D�_�5ݣ�8y>K�H�g�XZ�@�FH� O�#��ؚ��8��I�
l�C��������&��.��0d`fg���.T��d+��0�"�Ӿ|W���Ny&���t9������R�]�Ryb`�5��"j�n�>[w)��eo������~0^�[9��P�~{�O�sOKe-sT��X�M���ns��d��G��/I�ʎj���uDk��G�c]*�}T�0z�o� =bR�쓻TQ�LM۞�[�S��=a��H&��T}q� ���S
&3tG��w���8p/�*0�� �ߠE�<��ŕ�3#�DA��)}���t��B��7<��C�[��u��HIS�fR�$lpiVKx.xja�UZk��>�P�5�O[[��QKl�Vp,)�gr�گ�~�R������t�n��}uǹ�؝��ۦL�RZ��d��w���C�Ѫ�[�Rm��5�D�NP�J�X.�>�:q�0��4dx�/a��p>�(�{{.�Z6�u��Й{�����1Y��p+-���q�[sѳ夔��\�:^�W����V ���{���5B⺹鮽�Q��+��YMcN�Φ���B������wc�l�Ǆ�,���5n�&�n�=h
���L��v��;���>�
������K�~yfL�س�j���'�$�4����'�TK�-��*��5pǠ���u���p.�V���:�%O�ٷN�E��,�W
7u��xߪ�Wc*<�1�\R�y�y�B4�|5*W���ގ�5���Oi�.>���x��r���?X�)�V�E�Z��/�������(�Yƛ�� >��5E�W[XD/��6T��5����/���J@̔Ft��P9,�kpS��SR{0a68]��fȔ]*��5���A���k��f���'�l-�a�C�r� F$�	q���M�E���j�DI�-<]s���^�ϲi5rT_���0�?��j�� -����X�M:��2m\���S�>>��x�e��۔�ڬd��[���ta�!{I2G�]64�>iVa)X�,��Ƚb-$0����e*�
DL��(�����x�T?�TH!ohJ��f���r�2�=٥c��w�}n�n;��D�X�rU��5��ZCcx^�����И�gp��B`4.���+�f8��=�.N�oξ���Ido��G��S"E���L�I�9��`�_?.�~��CQ��9]
�RZ$"5pu%��f�Mـ�z���D��}��]��~��pY��,���<bS��J�J�f��	�7j)Z�(֌���J�W��=H��<hZ�y����3J,�I9"eK�c���=^�&ndvA|��f.T�d�J�mjc�3ԩ̉?��hK�3�h�́���YL���������/�ݹB�������[^t4+�":���I�n2B}:tp�+��B��m�K����#u8)�������]�L/��V.�y��:���;&��B���G4KSUCB��"��fH�b�T�uw�Q��y��6�Dp�`Y�
PT"���
��1�@��B@�a��� �4� 4~)�Y��co��v̚�l���#�'��R����I�E{K�!�||���W��sͷǢ�sv9hJ4f���}�� $��
�g��ǼtTK8�ʃ������D!rN*�d&e�؇��i9�GEw���9�RD2@�R�2��3%�����������O
�9a*Q�<��5En�qk�f ��ff��Kb���u�[��A�)(U�������A��qˬ0Q$L���;��M�g�-,is��cG�i��o�Q��b�mCGEn&����sBt�� &�`����³���% pB>Z�Vٗ�����?��V1u�WM��	ak���E��ۂl0op�7Lk�]K�t#�6�Ёd��vb��v`��|��D�������j���J!v ��Wڨck¯�����M%bF��p�/;i�!]�����p�y�j�=���M��n,d#N��r��S5�T�6�w���H`B��N\~�P3�-Q_�h�� ���O�+m5�.>�8]k�ױ��W(i�䬲�&�u��'�x�]UDw�"g�N�r�"���u�5�n�2��gMFt�"`}��~���`)X �[�C����	��kݮRA��6"�����a�k�Gp�/��)�2p�\cf���H�d�z+�؃��2�dGi��&(�8��B"©�$�UO���"�ƗyN�4_��lI�MC�z��=�J{l>_�6U�����pӀPBއ�
˗'t��M��7��w�pC<�-�q�g�H��zݵpH����=ZH�	��gb�h���O����N7bz�� 	��6��g�D}�u.����]�����5�ˏ	^+u2��8���3֩&>��>@���Pf����&��f�{�۔�,&��F'��r�-�7������������~�ݼJD�>2��~
�Rz(24MK���I�tM�+푌�z��/r�x�ec���,�3{q���8ÂJQ�	�(�)�W�N?$�@���ư9�����&�{�R��O�J�Gt|H�0U\~��%�[�M�g�K�W@5WU/�t����Y���_�?���ο����t��GN4b��ې�X.�|�8^����K=9����V���v��c��ħ�õߥ�	�e�6�8���%>�E�����CT${��������١g�+��~"�������`�W�<:ߚĶd|� �P9|sk��m�!�0k�]a_�$�4ҥԉ<j�������^Y�����؉}���wL�Pڭ���C/i&�:����!˚J��x�MVkv�>n��(�K&�&�7�U�;g���w�U\��R�jm#wNq�3kݒ����(&�,U��j��aL<����"F����&�'��H'����ۯ<ʙ�<8�W�  �m�a�D�r�J����c)$�i_��|�`"��ö(�!��$J[2pu玡{���|�����1{�L����TవM��u=\��q�[�E�K�l~��,�G�ȒHjET��w�N��KX�Q����g`�Ğ����p���(�q���;Q�w2��ry�U�p����gr��8���Sn���3@�5�����K�%<->2�,�C����o��\�P���*�P?�O���lݴ���z�$g��Z�5Ss��$qq�V,k�/��C������w�Ƀ�L�_+���5�腠�y���r�Rj4����Y݌I*�~��v�b����>n��UQ5�����d��&
l_Yu>�Ҵ��==�/?��;�RF�YsL�=�*+�fx��ܰr��uQ-���:�g��lV*��O2�����{�q^R�n��ᖗ�|@�ި���5�/ց ��F�#p{����3-��;�l��S�8uh��:�tk�����y�1ɓQB�%Ft�fA>�lz��n�#�u��:����EY�:�mK�^�L�"�+]o���Hװ�=+vgN�`[�<�Y�̗�[If�Du�lS-:�������#`��+�J$C��@Y�,��}EQ#
�D�$�2ϫ����l��0Os���TQ���I�!�#vc�X�M$!�.�q샞-]�ǲ��D�4?��dd�D:G��^&LgI���8i���45��̓ZgBa_]�6�$����ܙ��|���I��;�+�h�%���d�n��M��"{��4��~|O���S@A����\
�P���gƶ�,],@�A�5T�,����ۼ����:��~��z��+i+�L-dʊ�;KBٚ)��Y�ORMͬښ���N0�f���a���?���-���!,7Wܻ�u�5'���B���|���EXG~�(�y�VEP��t�U-���BF٬(�PM>S����|�:p�Xp�d�Ѡ�:8�˖��rN����F~t|Q���'G��"{�;�n��8�p���D�7!
��s������T�����]�f�`0� ����a��9����y��ҵ��͘UG��}b�=��_pܷ�����ּϿe�=ܼ^�IKN6ܠS�,�
���=Ð���2�~��3J�VB���:�_4�=�X'+E�%l
���@�5�i��M�E������lb ��^������H X��ҳ BpzKK_	]����K߲�����>��},������VW�a�EF-T��Nf��i+���'�	}�gK�������4�:�����W������� ���!�yqy�t+T�ĉ�/��R�YS�����[���������]��:� ����|<��(�w{h�_�TJ?���R��Dg�-F�p���A�@�
�u �i��C��x�	��RP���u��qfr����i��?���?v���SԎX�5��G��[)��r�����;?����3=��!��/[/�lf	O��u�3�2���8pET�7\�w{E�ps2 �i����Z��+2�y���8 �42 [�T�j�~'�]�ʿu�t}�]�\F�:M�9�'M����\^mL#�>�?�g�Sx+�Z�0���e����~bL�ѝ=�Ϊ�yEJoM.���"��h��\%�;@�_56Ah�Z����b��t����w�;����p�W�$�?`�b�a������"M�r�apZ���%���uJ�*	Y.�`����E'HIG��p�IŇBJ"��i���M�D���;��=!;�}cr�h��e�t	럍&=qR���4�)������[Qkl��p�=c�03s��j[� �j�+PaO�7���ɵ��Q��h�؞��y���i���{�y�e[w! D ]�|�pG�F귮��	��X����В�,����@��=��W���?]> e �ES'7O��
�_�Ր��s�fؤT��:n�~H��%�t݌%�DIbE2�!��(c����@��=����#&l���2)���:�(���2���ZC�����*2p��fa�=�U��f� M�W���������}_�$阭FP�Aa���;�җ��Բ��쬩$�1J�t�;D����;��H�v6�Hd��6�J�y�-��PR�`{�x��P�솻"�E�&�<��SO���Hq������@��"��gx����@�y��o]N���6PjB>��X�M�y@�*�S��~^�-_Oх�P�M�v^X�v�_(�J(T\)T��>�T�u��Ϋ�V�aK���!��[�*N�t�ւ}��q�K����k��=k�� ��&��P�&JoVD>�qf	��]h��~�옫&~?�T�/��[�a���h�_��<1�H�sұ��B
��.f7���(~�@C�`�*V��)�-c��է�"��pk"W��IEy՝K�b��`Q��V��hM��Kn2��'�����Q�j!2�9X��%B}I���mO|��N��8�c��X��J�0i�i0���Z��l�.Z�����v[����]��q��2Бp���=�ƱR|m���	լ.�-�W|��]ڵtw8�ܺ\S˃��^B��;���'F MY���.��KQs��?��y3�8Ӫ%��V&� T�I�����CE�u�9����\a��/��Μ��������2x�+�sz�ڀ2Z�F��b���ݱ�9����l�PO�Q�~Uvi&3�>FcPJ����A�i����!�\��(Z�e$#��B�����c|���Y��_��UQ��v�^�1}K?V���Lr O4M����J���`�^0����@}\�݀�rH�1��M67��e�쾰Hqd�Ye�Y���J�_��҇Z)��=at��bI�J��T�vٔ��ʪN�֚���^�+�w���/���=������wU��s�Ń Q��(��^ ��T��"�=��N�ME&��ҏ7��X^�rR|�Ц��������a�~d�X����>������m~��rm�ѧ�c��Z~
T6��R`i�zi���]�>6������ψ�a��X�u��$YI�@�V�@H
����/%�yڶ�Iַ1��z��`q��u��8a�w�f�- ��ӿ%g�(�=�m�������q���R�o��𬳎���W��A�t�r���t)��#�Ż��zWָ�zZ+a�Ru]PV¦�=˿�M4k�Nn�m1edj��g�2�����8��;1K(]y���3as��J�_Lȑ�"��[I$����,�*�. P�'ːxx��8's��Eb	9��a�Z����r�@�&p�uR/l%R���TB�	�NoA�L�}������s��`ኣ!��>�;Q�	o�tׄ����Τ��,-�pz��H���x��v ���:�Ƕ8?RB��\��m�:���̆,1F��b�?���JuG��3�"�
A��"�2�g9ܠCM�*i��)��`�U}��4�֧f��߷���Q��ߕfQ{�
.�K\��}��1�n��/EZq��\K;�K���t�2s�`��̔�^�I�&`��?�e���o�A��B�@|�O�K���� �*��r[C_ta
b���"�T����M[����\�V#�Mjݎr�{�8�qcZL�75��h]���$�g����� )ݵ�J_ov�u�X\��&K\�h�F�;k&�����E�cB��� �������v��_�|l���AROA����eR�����|�����H�M0 t��T�z"���g6��i��8����f��AB�|������4��ʾ�K�G|��_����'S�KϚ:�\�LN��#���r�6�ѽ��>�ڵ�oI� �"�s�#�bF-|����E�����{�$V ^���(>H�N��$��Itb�R���Mʄ[�G8�� ���
*x�@m����w3����ϭZ��VFE��Jy��o�0�`�۽�d�*7W�R���8�Ct����ȫ�>}�06[
P_�AҒ@t4Or��r�����A�-y�ѱݼa��~�_8��M��f���$�Р� xs��Mm��b�P���/��HdB2u��Re�:�yR2�+�~EO�J+�O(f+x�Ğ��!��%�1�A��0%�� %3 g-���T������~hS~����&�|�v箐�!�r^�����!d���u�@S�`��dU�0ZrU���.L"~�=��U��+��>g�N<e��1R��� ���,Tg�6��A�̲�ŵ�qhTC�k$r` F�Tr�V�_�$�}�Eߦ
�9��42��WY����+_�MXRS��;�$��*�@"g�axt`=��T�����:/��D/����*�l�K��؜�d�2�t�+E	R�g�E�����P�w��5�I=iT���p���C�l�\�tCY�M%�/g���u������/Q��]f*����5(z�8Xp Q,X��.A���Z9xA�w^|�ݦ���ù*��T��m�ӑ�/F�f�y�Ì9�7��t����Z��ʞ��	���[�FlUKE} U�p� �1�"��b)�A�@1��5��K���ǭZ����R6�s�;4�O��+��f�r`���L>D��֖�S�oi�����sէD"�[�ρz�QBA��2#��Y�r�2V�n�9Ӧp#�V2�E=N��'%��Z��)�n����1cX�jJ��E|���{f,ik��J<r�v��X�HF��}�D��$�<s��o�|?��,+
�ڭ���?F%Ň�*��A������` i�]O
3L�� �Mik�M������ݲ��X<�e1X^���ܣ@[�My/�K��3����m{! uv5���ApcC%����\	����������w� iHE��i|��	"Ɓ�0���'ˉC���T�	��z ��K�w� ��a_Xt�^�e�>shN6��ف@͂��v�N�a��|��>�X=٪�Q|2�E O�K��1�_������E�w*H-��D�.�>._��pk��He7���-�(���8�(�_f[��t�<L�a���J.�}��v>��y��|qK�n�gr�
����ߟ�W���/
.�=��-��E�t��x*��e�hg��	�(�	O�Ra����#��&1>M��O ������1��Z�����T�wd{�%kn��g��2�7�q�^_�UFy%�y[��o��DO;��sz��I�O�m�w�1a�r2e��E��z>7;q�
Z�y+��V4�J	H��'X�9%���Q֞q�y�|u�o������[ t�+&W9 0j�![�@C�_�t��9�ZJUx���طA�3�3�̇�}�>�L�U��8ޒ��4�>`��	�n]��~��Ծ����� ��)|ђ�5��GlB�~&pW��� ��}�8g��bg�7�%��N1�?�:R���E�rV^y>c �MC�&"I1��υ�e�ە� ��SL$�}��j��cU����+JxaϞx�K�?}}�54��y�H��x,�vX�n����׍��՚vڃ<����w�ա*9���E]8=�Y�gs$�{%<"4�,�?s
�%��5����4�Ŕ���P�3�X(5�,�(��ƴ�5����.Ep����H��P9�����sЈg�WOR
n�]�sONM,ݬq<�/�9�J-�a�ps�����3˹��M��Sy;U r�W�ٝ}��Ë������1u�Q��Y �~/��[�n��,ꃋR�0YB������(�τC/ӭJ5�/�K���TISf��-A����;q�,I���t�3����vl��d�g�p�H*Ni���N'׮	63_����r��c�;8�/�0	�f�t�~h�ݴ�c/�7�I
�FgQ�!eԃm��F�J5���{
�r�����eqSU\���I��!qi0�
�R��#�>Fd�-ez﯌>�q��#\p)1a�Z~Ɗ��2�YQ9��1 4`�V-�;-$������r���"^�~����� +��:~)&�����02�
�4���V#^0��m"�Vםx��D�)�2$L��`�����OH! �C1v����<��;�䠏���u_mZUϖ���v�lz�
�K��r�|�^m�]��o�Ǔ��x�&w���V��"6j�E�p��}�0v���"��S[��;��q5�4��1X����4�l�T_]��.ن{"+n��6��qVHȭgW~��|��NI�%$���0�+�Y�>�@�����¯|{/-I��ċ�����"��'�7���`vJ���%*��{%8
�уZ����v$2��x{��Ţ	C	'�Tcj���+)������g+X���kzc6:g��K��ލewQ��&`z�M�P�_�٭�I:�hY�ecڎ�9k�H5�I>u�yb�����^� �� �]��� �x�;%v�����8L�d��f7|��}]U���.�+�������8�r� ����=�P0�7C�h��U� �I�	rr�3!W;캒��pu��߂�.�"p��[Tnq:��Œ��S���tc����gS�^�D��p8D֏*^��	�{����N�8��Φ�:9E�q�2��BV�x(=|A!�b�w���^�4y�Y�SaS��v&[	��Ή9�q@X�8�ΌMv5�;8���G�,h�䊣AEps�gZ.H�:N8*TcʬZx>|��Y����Kxʫ���pBa~@<X����|���'#��S�}���w[�T`<>���bK�F*�_,^�w�Y��C0�G<�yr�8�YaƢeu]�Z������|�[�r"B��Xr�r`z~&唫ާX9�Ăz�p���f���e�e�]&ց��	'v�lŐ���/���[���/��S�fUQ�NJ�Z|SA�5X(�qX_x�wt�"`�Q�M�v9�7�/.�}����-��l-����6����Q�C�� W�af����#�}���옠Q��{'6�a T�P�'�s�u��/^�m�}\�p�^j}���ܾO_DtuSI'�C���P �8��8����v���B>*ո�I95���]���b��s��U�7k�*��*:��uT4Ά�{�n(i�����I��o���ݛkN&��Q�"�P㮇�`�9xۧ�U:�*8�%�4a����5mw���{-X������U�
�zA
�zש=4����(��o�\=��@�>� =�a�^�ய��n�T����B�[z�OrtK�9�To�N�b?��]\�c+��-��.��+�p4-��o����(��żz"��2q�9������i�T�\7�x6������>���v�Ǫ�qO`K�2��,H,��Z�B$Y�wdW��F<(tW���E��r�n��uAz���#����>�[Q��H�����H.��Y~��I?�{����*㼁5p� ��1�\�f���z��
~P+���7�\�� ���D���J�Q+�_�@mR)\�!��l���)0��)͊?��:�$t��$�y�+���G@�O��vzl����K��x�>��L�c�(,��£��lǂ��R4Rd����yѤR�œ��O=��^	�_�9J$��� ��~t����5۷7JKSb�U�)�U�������&�tj,�ltѨ��	SR��NR��&��e�z. rJ~}�O��kZ ";6����!��iH���� o$��"��j���# �Yi�7���K%)BA��|4�"�Aғ��M`#xD��}�|�<3 r�
f҄)�L��5M��bjB��ow��j5�C�Aߐ[]`�>lf�
��:DD����ߖ3�n����G, ��V����^�8������i�|+�F�3gKrA0��A��� ����\K@�V����/��՗���Ո��me�|Sgy������g��Qr�ƞ�e�#/���V���D]�=��u�cS�F��Q��U�
�H�<���ʉ�#����gS�����p�=����'�Ǹ~�����"�K�el؛K�����Ťa±r��-�����y7�[1˩�����)Tw����}v=�"�0�N���վ�ޓ�dL�W4��iKޔv+Ĩ��$��;�?�3��bDcu���Z����@�+-��M�{���L�Y�^ 8����ϙ�Z	�kv!�i��h7Pb��f�c�5K�R|�`]V��٨}��;�� �J�r����=)�=�Qe���%���1CH���B E���Ӥ'��y8�Ԡ��kPG]���d�r��(;�#�{�?{G儦������bp�@��iSG7'h %�O������_^\i��׾�Q��+��>�T����C��;�K��*Ԫ�q}D=����qn�NOxHR͆��7Q�Bx���B!��S��,�{d�F���B+y	�����T��e���%]k�c���E��;�	�K���s3i>9�>����\8;�%�F�W��e5�����>r]@��ݧ�1 ,΃�#O^R����R�����+I���6���oGIz!��y8{V�5��eS�Q��,
���G�i���T�Ф�d6�]��=Ͽ㯁Z �S4��2U�++�/8�"�F��^ͤ�v���H"wf����ڊG�R��4
}(������#Ղ�����+b4A�-�����&��ջ[�tNl������з��Sa?/<��ܘ�:�WV7��Z��FmAI	A��y�ޕ�,����b1頯�[�y���\�40}Rb�ms=&Nj�d`J8�gҰ�%�A�K�n7K8��o0��T8�M��8�)��*��}��wħ�9��Ѕ��s�A�Q�5��ọ*�y�|ŷ���ރH�����˗�R���CGF�9��7�'�b��������OW��z��(�S��FȬ��P�B��\�F��O��PW�<+�T�5�%:� U�[(�䣞;?�����Z1
�y���=!B�P�н��{�>�Ww[Kx76��x#��_�c��B��-���p�F���3���������ݷ�6C��A�bacG3����Iܐ��AW��T��x6�TcWn��G�0N��g3�K�u�\�I�;q���.n���s]4ᢟ��:A��&b�~�p��Y�Q�(�\��JXr��=��Ifv�zn��D�z4w�p�1��0,�4����ӥ�o�W��~е�F�#d�8�,��
z��ց潤X���"@VY�����z/�����!��q�Pj�Qۡ�fG�<H	��w���$N��̫��q$U)���J�=<�O~���y�h�?]ڒ�j�����麌8þ�x��_j3:nq��6��T�$ŵ�<<"�6H"�rƬ�������5�N�z�GEt�z��2�۶I�5���r��R?�JfzHPD�}��/�W���W��w���ή'�RW�
��U�5e���v�qѓL�h3�H_3�8q.1�ڝ�%����R�WsU=Joֹ�\�-�.p"��Q@�h��j�;�C��o�Qb�y���u3taz�@X׎�_�a0�9�}P���ka��}A���Fm\�[�	L5w\OnA�q��<4�i)�w��8�����)�T1>�QX�у�#<z���?��Sy8�� ��3�[Ъ���ƫ7 q7ML-��7��.Q��s#tZ�EhV�a���0k��xQ�"��L�DJث����)z�V=tWUD"�R25*�Ã5�3ޏm�d:��n.�e���+�I�������n����M���g&�rzk�A
�x��A�P5~��1�!(mmr.��@D:��<���>�A�uG��g�O*W.�`�p\�j��~ώ���\6��GB3�85`W�C�f��zh���H��<u}B�aϕLU?�eWd�=��Mp������Т		��7��A�l�	æ/V�|�=�R��2��l��J�`���8c��'�}n)��!+$VB�� &}�t>�m����ëɟ2Ȭ��
>�`�e�Y�=5�3�:�*��c?��x�V����䄅�ˊl$��t���%4ķ�x�)����6Z�y�ή����&}I��AK����.%̯�T������Ws!���yO��	ڕ�y�*sw�|H��E��Y��Cd�D5��ɳ�$�Ҝ����s`u�r��R����	�L����q�Κ��	��uʨ~3������A�4�2����`�*��w�O��L *��5w[��T`P�����>��&��
u])�Z�N��N��iux�u��z��z�Њ��H���>[ܭ�<J+H�dV�9�Q^ Ώ��t<�]F:��F�������8�!�NG��\S���/����A��Pq�#�g���Eȍ�n|��1�BN�	(P$v���O���������͐�?0���4�&�c흘��]��������*g������ݧ^�_���n�b$�m�l�u�f��䘜��=a�@V�y� _R��n�2WGd�~��Ael�*���05u��5@oIv��6`��ޯ�쮛�f��4R�hmS��d�Y���7K��q����
ے��Ĉ~���L4�J�g��/��u����Ť�j��kd�@�I1�3��`.^fï�;��p C��'M'i�f �L�j{�$:�Q�d6�5�B�3Ұ٧OP���	��3�j,� �TU�%�	`����@wLK����1 �ܻ�/�ɝX�jV<t��)Cfd���� �W6����j?���`ꦘ{00ؾe�9��_")���'��P����6�"ćQ��섴"��9Mc5���1����fm��F��a���Rz��<��{��a��u�;��z��a1�
�����ێ�Z'i�)/��#�*@��Ҋ���
*OK�r�o��!r���#"o��c��̶��E��[���掀;�������T�O v��R4^�/�9Q�ǎ�-�v��]��45��<W";e�ߵCP�4]���i+����U���jh98�wN�/���b�l1�p���Hw��h�Q+�袈ζ,^�g����5 ��őWK����0��WJ����#�a���o��ICi�� j��*j�VZ|�������?��]��${�w�WZl�t/MHb_.���(O���g�J$Ӟ�(�`��%<�������o��*��׌���	zv�Nct���fr������(��˂0zQ�y��AkR����ck������^�~�m5ib�g��.]8��rY3��kn5����D��{-�}x�mv�9l?�����L7���"��`#ئ��w#��Gxd.stt2��^�6� ����\���\����\����L��c�׷Z��6�>hs��<w :��ю��b��ŀ�/����R����C�Q�l���ɹ��@@s)+�)T�P�������%�m0�bz볓�jͥņ���,W�š���,	 �}��x۽����B0w-������n(�w$Ĕ��KT<��	Ʋ�9�SrW���h�!�$հr����\$�G�gןK`�E!*�d���)���@J�r�B«��צo�i� Pd�
%[CƸ�=�i4��6�-��P5ҩ]�*:�n�k�N�J����|����/��t�p�.�P�K�-C�����B�p��d0ƈ�����nFl/ c��)�(���.�nyڒ���8���	���'���z*�
̆ǷKŷ�}A���7�5
�B�{2uG Ł��[�qh�]d���R�Ca~����[1��	���~�y�XJ��ٕ>5m�\���S�2䃂O ���v�SQѿ�_�f�7�z]��\魾[�|v#/)��gCg���Ҿ��֌{�Cb�̔eXw�7ӐT/�S��p�N� 9���	Q��#X#��-��Qo��{�~�(0FY������̝㲮���l'Y�K�>O�+�2�״�Wv�$���hI�HN^+�Ez⨝�d1LT�0\���q'Q�+�E �Բj�IP���C��Oտ�X)��8Vqx)�ZR��D��ׇ)]���ޓ@w��c�9�k<�W]e����f��޻����X�x`��� �֐݃2��f�J�H�o+_э�An���}�H������@��oj#m#�g���|$�m|�8�-��9A�jDNy#�OihF�I�$hu( �JO�B�Ii���y,%g��#1G��<":�L#?Y%��Fͳ��~6#��Q�!�I���V�6��B��r�"��ڎZ_ý���3>���G#�ӡ�q�9G� *�ww�/�#x��#���)
C���A}4Jw�o	S��O2�,c���A ���y=7D�4ؖ�М��Rf	{��XUL�������2۸�v	�,��Y��벓��>���/	�򚬓�Y�ń1��/�Loʀ�T�rO0t)uU 9ԮƓ0G�����0�z�-�_'�>�#F��(&թ4���Fu�H(�0fm��4����Y�~�@�8ڻ.ʁw�)F�oE���_��\�|3�˝�O�����l�H�xC�yv�W��T^`Lu����ݧI�Qj��D
�	�X>��@�թ~�-Q�t�6 #e�6D�l#��`0qS��c]���u�xM%�kB	�!TkU������\X[uM�D^m�A�B�2����-�$L����I� 9{蔖жC��^L��X���`�9�rlSs���u�N}�H2U��FT ��m�R��BQ��P c#���>��͔+9�M��ڈ�SGY���y�	Ԯ�M��X�� ��d��I���̌�k��)]��eӤW��\��,��X�S�	�8\���騘���i�� "������f�z��� �ƌhc��j�
9�,�A�-��B!Z����W7��^p8��â��e�F�Bs/(�v��"�-�N.`\��|%>L����97Gc�Y!�F�.1�
]��U��<�[%�tOC�� ��/��rVGˆ��Gϭ*}��s	�U���'3���1�#F�E�@�����S��x<��}mh��lّ�O���1�m��'��y��B��M�j���/W`��,�&�����A���x�D"�£����қj�E��]q�IF)�T�cZ�q�Z�ا?�i��Y�!�k��75ά�÷߰�����pFuMQ�r�k|�r;ˋy�ڥ���{�Qˠ/�#}�i�e���)�#�]�`���nZC�ck���'?F5����!j �EU�����%o�!W!za:+J���k|c����3�wج�9��tW�,K�R_X�����,�	Co)RS�s���544�3D����	�	�؈#��S%����]�`N. 5�}���^�Y/��ǫ@U��~�cD��W� Ix	(�E��3U���I(�nx	@6�DEq)ε_��������z��	-�J�|�c ��C ���V��jb����g(_�,�t�^a�@xI���d�Œ�ų�z�SD���*�ьd�XQ�k�%��F/��on2y���0�G/B;M��)K�ӎ��ߨ�͙E�h�c�W�f�#�#1|&V� �2���2��B���G���q�������޳I�hŘѫ�=��$�x?�%9�ɺ.٘U"�V۞����e��*���Y���V� �t��m-�.���|�O��L�����!2ۊsf�j%�����m�gz1GL8T�y/.�@�,��@!8�[�ï�S,�����PcB�>8�g�]�H��#�#g|Y�
_ݱ�x�h<r�ѧt1�0R�@g����؆�"�G<��r�����'7n�~��X����s�Kv���ܥ6�~W�a���g�pÈb[h��X��<C������X�)h�������8鉣��I�N�K�����K颓��c�*�H�q�DSp0����k����
�r����M�ȭ�ν&�Pt�t}�O��Ȧ	YL#�g.!*�P���>��J�m��36f閊�75�\� ��|y@N��z�\�q��e#�U3�S>���+�2Y��=��ʍ�Y���a�-�ĸ�q6��{���[q<Z�p�\��U���Ar�������jc�c���awSc\��	gun��������ke9�`f�q.xMK�ͽ�k�p솔�RX�����
��MZX��l�Jx5Z�]��^)�}E��3�fjq��e{l㪲^m���Ml�7 ]��JgYWsMy��o�ϫ~�
�����#���tx�&���lR���ym�W�qq�.4(Qt�;��@p����X_���5 �4D^�t���:CϚR��_nu̡�uպ�"�n+����~��� d�;#mv����o�r�6���/9�T�(��5�JC���H�8dX�_�ᅑ��W=�B8ߋ$�d�K�ƈ^�N�9C�C��@��W0��+A5����$s�����@U5���k|��z�	�"Ms�z�0j�#M�Q'șo���[�Ɍ>��3F��pw����
�;܆��6! �0;IK:$��i7p�����x"�3�j��j{7��
bؗpq��J���NG�ЩQq�%1�*6�1YP��g��'��v*�4祝�|j`���л���v8u��^+_	Hף2�]��0}��j�{X�ap^!���$�\��I�Y󤣥���[X�J�zɼ^8�$�)5w{�^b��O)�`�;-;��� 22�u^��f�l�r9�0�
c.&�C�;�~��0�J����{�^yH�G�:�����k��N�p|3ײ�qm�t�����ՏV�7i8q	c^�1��N�CY���-�*^�{E`!��a��Ny�5|���6r�Ǥ�� �(3R���/�@�M� g�O��UKJ�3�̘�1DC�T��Zg@�xsEp߬����	�����>�ɸ�N�dS�ӹM�S̤i��"7�E'�{��a���b��a��&����?h����B�}�2������T)p�k����Aw��\�lFW��r�C�/�3}�)//'�\��L/���W5D��(�'߉��~�U�"1�Y�^�����b{��?KQ���������R=�ѫ�t���H�Wc߅�~+��Ź�
p�jZGJ�:�j�=�(P$��G����2�,�ԛ:�
�@`��C�,��P�Е��EaoK~k�#���E���E��=��l��ꔩ$a� ����� �UC&���J7��;�w���kx�mܗ������oD+�rt���!���'>����M�"
BO����HX��P��i���7���M �r<�%�Ȓ��`- ������H�"��H�b�0���0	�q�顚Y�چu��5�g�ȝA�Y��F'����[��v�}��J�"[�n��|u{F1��2|�n���un6��e){j����C��S�T��tw���	��Hj{\2i#K�)�?�5��n[B&�T�� @�ƙ�1Nto�F��mw�[(������A�L�\����Ro��*�,�ԣv~� �g��P_Z� ��|�T�U�%?Gנ��73z��b��c�e��9�kG�ҵ���k�$������-r`���/�	=;�3����o�5�qL*�G�Y���{<�r[H�������䄡�S<�QҩIY*yiI?���Lb)��:�3����_�g\�e�Bt����ݛ��`s� �����������:�U>q����~,I���u�5i�Lp�Z�V�ԙYU��9빕�t�A�*�cIt<\�̰y=�Do��ڵ��������UW-<H���[���.�5P���}X�K��a���P:�#��|Qn]W�J�3eN��2H�i}�H��a�<��Lk�99����C;G��pT²,qr������(���� �cˀ�Fbn���%4��~}���Ć"�iwm�3_�Df��#B��T|�?e��1ƙ��~#,���ڑ��P�v���u{SG�f��`�BEq��WFL�|�e{1z�ݟÜ��£BqT�B�M�ç��8�'�	� 1����q't�0$�S���<�t� �l�)�70��B��]���-���H�!kl��˼?jj���:F�IK(Y;ݾfi����۝Zᰧҿ]�zlZ͒5�J\�I��F'}m��N�h �Q1���e�e������(�_eXڹ�f��G��qf�W�[5t�vD�9�*U@mT<�:���L��ہ�f�N_��(�Rq���J��|�M,�P=�p��O`��b�Ar�#M_��m5��T:7gv&���G���z�:�=JWǖsέ�ZM��s|�98��`�B����Z���̆�g�ک�����h/�(��A��#�[�����{��NYD��vp��;�2y[JO�k����d���&��VS��ܜV�qr�e!���2�o�3�as�w��Ɏ��Y7�zwGu��wZ���V�23�����행�����Wg��=��-��������N�H��!&/v���s���p$�fϜ���IK[��"g/Xx�h�3&�1F+;6�o%>@{�Q���uK�9V��֪���;Ɏ��1���p<�E�B֗���kd��<~�%��N�Ѝ�]�e#�f?�J0��z59�3'�*�p�2�k��
Ns��ja�}oY�!Dq�>6��7���<���.��y���Sy�,oڧZbW�*���j�Gl�h<��f���6��\ n:�gԿ�L8��;�Ϋ/��kT&DL��^��H+k�	�7�*���t	�bdtN��V���lAC�(��э�.qjM����"(�yb�yE�[����i�H��X��>��=��B����9�y[R|@���dr5�hU�{��%�K.�R8���ࣳ��X*u
u���ֲ�H'Pnp��b������� F�0 �c�jbZ(�|�N���wJI����ۻ�I]�G �.d�ȟ��p��i�r8m��]K�_���{�z��0�Fp���m[L�$�!�hq��1���2U��ġ�b��g�`�Dql��WA�v��Ekp�Tv���(�@�����!lF!ʎXC	���$�}$^��b�$�g��>�pR��R�6����
�5� '�>]?9���YB��B���)��:Yg�@n�t�H�)`�}�c�����Iv=Sd]�"c'chԪ�J�ؙȕ}�-��\�
rF���h�*������v�(�/pV��$r,F��.�[k� Ȅ��	�凚Љ��W�"��5�9o�'�nR�<v�cN9?�!�Gs�*UǇ�}4��I�r���zS�tл�^ ~[�?��5b��YlW��6_�q�C4�xr��5M��;BN	�����_���@�+���̞\8%��ܑ���}`kK}�ϙ�Id|q�M���)��@{���?��Ày4q�ŝi5�ԇs4�Elm�fW~��-�D����TDa��/K�O7"�!��Ļ&+P�r��9U�.�[ĺ�ͧ�� �2/����rjx���wh�D���&ys4�/?&im(�"|���W��-���JT�����76r\?��o��f��s[���>�p��3����w��cs�)Y.�m��@���I���xY������>� �Q��
�E^�k��/-~��r�9��W���H���)x߳A P�����N��o�6�JN' �|M|��%r����� �T�t3�s����=-�YO����m��@]�A!��͖�����x<�{]⢱04����b˔���7��^�SIv���3�Kr6ep�>1f�'�3/�M@��<���2&�>(�n�N�/j�U>Ǎ�� N*����N<����W��7om��v=�{�[�:���� 75�Ƴ����S����64� ǀjo,I�7m���-5�wW��Pa�ܢ��m��㏞|�oh:�S����C� :!h}49���Z��~�<�r��Wy�.hY/[~_PE8�L�H�x|?,�>�RG_���� q._7����[�lzc�:��
v�
\ʎ�m+h�WzZ���>2YR	 �9�\)�i�೽���I����7��+���Z�����"! ]Hy���#�(��ۯrI��Κ����޵D．rݩ����fT甈`��pr���V������|y)���枣U��a엑�։�<�v�'�Ŷ�앢M)���0!�@��G�@j�=�7��1��l%J1�n�yX ���}��7���!_�0ET�}�>N�/��K��<�Z�`���LX
�aa��$���j�=$��q��OgO`)}=��;�^.;�Tͯ��e�Ħ�z"l�n*���l�}�sH]��w���D�O�5&ŀ������b�4X��-���nG���l����z(��iq�� �ү���z {P����O���JDT�C#|� �� �uY\�nO��Ȃ�FF�]�����B��"����qK��ՆP悭�ma��l�I��9~6�����X����ja��v
��O#�HE��$�mr�
�|�����,�"���@:������:��&U���`��t1���p*���Z���Ppr�!�f��U#�w|��� ������|���"�$�M���qo�@��9I
#Ыl�gJ�OfO=��9�O�����X6J�F~���*=GS����aS�\�C~	C3�Y�*��,Gϋ�jc�����Ao�K[��d��������1"!���� �{+`Th��,�\M�2��K���#,�q@�X�7~̕�-�[���
C��#���g4ݧ#F<D�Z>��(|/���3=D��v�H����ռ7\
��	���0¹�BM�
���I�K�����U[�k'�R0b��쐇�����26�p��l�)��~���$9�B�B��.�B�Xp%��)�-�75�S�ARzwޮ�ֻ��Yz�i��f����LG�W?fG���w�Pw�y�x�f�$��+t�����-`"d�%7�{ls�\���
��m]_��9�~))a�ȟ�xm֛0H�#JS4��1%T��L��S7/����ha�71_^s���P����K��%�/NB��ȧ�����W�P�m'��ˡ�?�����6h\O��x4ȇa�4�Z�)�n#W)`�����T�H���i�(M��a�ް�|�搸$Cb���P,�;�L��^��� ���=+��T9����#�����#��<�8=�`/fYF������ 	]��Gж��3c��G@L�|8GT�$-�na�g��xjX�\ˆ:�["NG���M?H�^�����):"P{�������,cgNx��52�쥂��'{�
<:���It,	?�t��Z�A�K�:WC�Z�z��,?U�D��IE9y󹑯�|�ͼ>���;Ӵn���G���54W� �"�H�X�p�����>tK�Г{���k<�j%
��=�%.��6�*��
<0&!�׀$�TM��J?8���n�z+��d �5JH�k}��22a��THR�V��BJp&�;t�DI2)S�m��D!��;ʴ�$��*�SP3��I��cy9�3�%B�����b���L���OK<�6�jU��nj�8�H�� 䜞�|0�i�%�&]ʖ��劇�~Ô���N��Y��=�*C��գ{b
O�)����;�y+0��B�K�d�J��lq�d�R�}	�I�{�47t�j>�w�(5{����ᱩ��X���k��K �Kx�S9�( _cbc�/�Q�m���b|��ޯT<��b�'�8�u��ԤC�����`����Y���^>d|i�-*�Y���·�h�/���^���u�*"k�K�;��X��J�5HD��N���27�*��W�{M�#g[���i}J�wWY���mH�=im�M�-�������ȁ�..���oHF�h׮h%Ԁ�l&��S���G$�=��y�.�z{����� 黂.�r&3Tc�:D45�h5���'�M�_.d���<�_?E�F"��rz���6���:��+f�&Ei\�U��F���2I=�Хl6b���xi����Zܻ��y�Z�_X�/j��NW��C�J���{$�k� �
� ��Kc�K�/�-QC������!H��.�e����?�3�u����K,�^`�K����}M�.�����hiy�Ly-��;��]��'���	r�-�!��o�n�K��L��wBv��-c9g�ź�͡\�f��U1>��#�K�z�?�[�����R͑��4���>?��8�	�N��>���4��
���dVA;�԰hu���l�X���dJ����d1_�������� �އ��M��%�=��]do´v��L��݌;�1z��B��=�(L������vI��\dC�y��Oh�4����cO���B�֊��[�H���F'��1Y��F�$)ؔT!�4.���Cj_�m�Yj�i�V,�|li(C*����a�1��ƖPT�qy�T "(�������d�$�<MC[��<1�����L�� ��z��%#ҷ=N���b5\?iӘ��ǐ�4Zg��sB��z�E.�;��	V4-�]�+�!�xUЫ܎ڹ1��,���T���P�riS��LT����S ^���g}{��4�(�#̖���m�M���C��p�/�
U+���jO<4ᕓ�Pwe7}YF+��P�h����z��L�
�,��$�ר{pP�J��{�$� *q��hXoY��멶���.|٠!�G���ǂ.p|_��5�D1!M[�(���S>�<����l���iB������2B3M@������A��̪k��>6��ۨƖ�&��Wu��jB4��6��vԧ��;ZO�JlG|�-g���)?�tQV���G{P�2>�&9�mj/pg,�9$}��g�`lG���m ?a�ѣ ��/���O�޾]��j<��]��£�3�B�J�I���$2����,��d��40�x��%Vj,i�T���z05��}�hź6��}{��O~<Q�_qً�Dp��7>^�%�*Sd�i��[���J3���l�TXT�����묨�/�[�É�q~��NQ�c�L�O�:������.�UD����m�S�H��w�]�q�ß���(�7o����u��N�>y_q�E��~�R��c�A+�X�ǟQ��~��IUD�q$�6&���W�q�l{�����.��|���%�A�5Pzټ�✄�Y�����(-�	"~��e)��?�g�!�s>G�M�0�M�eb�]���R?h9�T�O4K�%LN�uX �v�\�Ĳ���{��I\�c5�~�	~`p����:�1wi�A�,��Q)������c�z�%�ް�.�����6�љ�K�6�R�H�s����>T��P����8�z�����XhFQ��}��/r�p.��b�gy��4Go���rp}��W�j�y�G
�����\?����"���ouU���>e�,���y��!a�?^�0ݼ5�|WN#�Ye�޼ \�@Q@��d*�4 k�Lm5t����� �dP�kz�d�6w{zR��@�xR6)�E�B|�e����3]��,x_s���ڈh��}roδ��#ð�*=p�R���;����/m��(�J��6�ݘ��D��+�5]ev��N�W'�j�"�軺��j'FKM��6�3�IN?�f��������:"!9���(��^&����)�5��2l-B�JH}p<ƶ�y����%*�Os��������N�:6��BlSO���vj<A��9E��3�ލ"���2S'&���磻����0��� e!q8	���G�[	DI���P*p��T�դ��<]�*=�Mᓏ>������dhG��z`�ԓ-�(ͻ�r���P ��Y���ut����i��7�1�<�Zbx:~^B�3�P�K��������9~w��lk�ս �&�-v�2��ueL&�V�:����ҰZ�T�$�����6�k���nz�u�=I�W`�^-J�P=�t f�	�us����+L��4K�3�f����r�L�[�ad�������(ک�+�����a<��ڊk?�n|�& H7��(��JEX�c�E5m-�ρ��N	m��'����dm8��6�d^��|/�`��-�5Wg�K���t���/��"힉�7�ފHV�~������1����ň��"��0��g���5Ro��}+������6�zu�hȬ�c�|��m<�&������Ԙ�	������f��EP<�҅p��e%)��GҘ��x7��9�
���=�����4;�3>!jZ�pNtfŹ��@TD�O7p,s�L�B���dl|�@3��SE��JNx1tTG���6ctg&��� ����Wt�A�Q��d*�uf���0/���<G�`�����T�����p�"�N�v�����m�|�䮥�:Z�"b���˞���J�����v'�ĺ��#<Z�/�	��^5q:q�p��;���]�F���r;�h�����؏����U��Ɖ��.͜9W�K�(��'3����}���N�6#SY��@f�����}�H�xB!A�8���)0��GYN�D$Xʝ.H��{G� ;��`�i���`0��f�G�p���s���ae��^��m��Dnd�9��/ذ{�ޏh6Ƅ���`*J�Wj�=�|�'k˶ �}�K���&����m30|�A���5�H��T�G���N�6�y�u��4�����U���8Z3V����S�{V2��A�j�ԫ�pn�/!�{_���V�_sGд!�ُ��b�d��E/��H⇫��G��ّ�<[�U�眲k��z�i���Gq�h	��ъ���ߜR�r(���Jnԣ��nՑ�MT��U�M) �{	<��±:�h�����Da��;Fj�8ʅ��g\k�
�غ[y/��۹����b�l,�.�F�"ijU���6l�l9b��`��ӕ��𷤎0�%����*�E��g ��R=�����Ő�R�\����E[9FGi��[�1��#$�8�c�0�]��VBi�oRN�ͅ�ky3��A��o��>���bA�J������i���5�ₓLG��IZdv#�mf��N2���X7��PE�W�P�F-��V�r_�[���x%�l�h�`?U
�w$�2	�3xu�;��؝��_d7�r{�9k,��M���F��Ծ\v�ඏ��K���G=�EZOe[��W("�>b2����Ȁ���0#֊
�S�v�t+�wMyF���h��	_�]TX;�23��pr���(>Q�6CQ��y��9�k%��B�_�I���H����WCH2�O&`�=2��oPRׁHs?C�o��F>���2�_mkoV����۴%Jm�j@�T��^�Х�R��y�!�q�E|p1P�~ءM&��h�R	T4w�4��0���bӁ�d�V��a�aB����}�s�j� ҳ��X�ߺ�Y���Wy�i�i�w��t���N�d����P���0sw�/����"�5d�y�;i�s��3����q.��k|;��:A��Q�{W/�z��)��$@+����6q�~����J�k��Iڂ�&?�N%S�rZ�A��T��.蒏�׏&�}�b�q�N�3���aԿ�4`h�7'R�hm��l�tȲȑ��f4���a�ޮ!���
��%�1�Ñ��Y6YyN��f<E���
^�����.�k�����r���{g$@K�����H�'cNQ�*.���N���^L�(C2Kh��D븸Jr��<t�O��R��sx''�K�I��yz ����l��Nb����
�C�jU���cDu�Sɿ����Z��4�,,��]<
a}�:Ut�)�^}8\��#7��
9����3��ھ�qS�#\��A&(3>a��g�-�p@S��C�cH#��~!���eC�4�E��=Tʇm���TGɓ�p���$�i=�����ѻ��*��1ҩc��t �A7��:�\��+ ��Éh>��8[�7�m�O�t�R櫎;!�|ER��b������`�M)��E�	B �XL%��)J(����ID���I�{څ���s>�y�%e`�v.�}=1Ȑ�������SS�,5��#j�R.�t~��F4�;��ј�(�O�X����z�P�܊N��+�4\y���x.�B��_yY�ݥ���T4~X�E*����t#M}���F�N_�[?�2^�$�T�I3@$,��(��I��)�b+�&F��=Q�*�X}���Dd���"��<���o4[��U�ǵywf&и_�Vo��R�?��s�k��//�1��&`�k�=,8R'5�	��=(��IkWwS]����?iDc��~��@cJ}"q����H�፹S(7�d ����j�t��g�NxO��,�g��Y`.��	�^$�+7�Z��t�b��>G����ڏo�}ä4I�=�/�[�D����&���5[7��ӟ��P]d��f�gd=s��`\�ˡ��%�������a��G�n2'��:�4+�
C�{EE�dO�*g-�_���GAF]�[�e��I ���{7��)�|Y��� ޣG_t+��
�� �����a����*�JS�)�ﴋҝ>F:$�����^5q�e^�n
X�:��29��5H���M
㧾]��6�(���C��_�`>��><�6ysD �e�j�!��t���_★t�d2\���l�H*fI �9�E�M��mT���iF~<�Y�Iv�1��go��E�9��(O���� ����v�FV��s�0J�$_Gtl~�L�j��|�о��<=��3�����L��j��8�����Eÿ�D[�Ȋ{jCX�+�	���V��/�g����GPU�hL��E;�{o5%*�u=I7�y���[�Ѡ6���t�B���9�Yp	��ՏZ�:�
��0+��������7����L�.˃���[+�	��z[B�wߢyE��O���k�����Z��2�?���Nym_о{x�"����VX�	�<��q�,��2��TؕV���2b�H@*�YS���%�	@p|�� ʾ�Gc�'b�2ۊ�^��h�D9�v��q�.Q��l.
Z+21  ��p��,�Q�u.I>�fj���z�D���"��U���S�\�c�3K~h�k$��0B�΁��
^�(���\��G��7��H�� .����f�DPa̡m��t�z�c�h[z�MFoC=�@�_cX�玤O��>�2j�vj�@�w�-��s�� ���E|Q�G|���_�i�:�����АMb�N�T�>����ҝ_G�� ^bzk�=٫9�c��lg%���������ʼb��"�����~��Ǚ_��g�(2.�`M�ڐy��B&�Sq���[�`��a�ڈx��>�A��+��z�9q9M�$�F�C�38$�fm0����u'�0��6LA�T!����a�uиI�U<F!+�-�z�B��^/���_�����ɈHv/�m`K4������F�	D��.)�h�'���m%u �2*)r�¤��?��+[�8��z�I[! ��*�$�3�w�[�+��A.g��F� jcx+�7��~8;BP�׾�4e��Mk�q�K�0�Y���&��( (s��d\���r)R�CwLN)A���|j�p�+N����+���^��L@���(��Z��8}�o�="��������#U[��_��CY�L ���/#ߜ������EF��>p�}H���;l���8p\R]�Q���Y��*'5�%؜K�*����Ħ��&}�p���?_Zڦ�������
iBԫ^MЅ�����-�o!&̟�'HG;�`9�PQ�c7�U��v:]��u�\o�ԝq����?�aZ�v�W��a�ت�=6S�u�z {G�K���u�K�Ⰽ�y������@$���}��ݓ�y�Wa]�a�'���h6�|�5b;�p�}B�E��$x�Dq��L�@���*f�����C��� �lx���DS�����kA����0/[EeY�?U���M�U���c��+�A)8�+d�O��;l�N����#�?���-�=nRz���򚚀�!�wrR�r�����}~�k78���9�|�H{��[�!���-2�u݈&���и�FS�ʻRo6jH,����)ф}:m����������,���*V^�+�`qx�ػ
��Q,��� W�*$�T8t�Mǻ(Z�*yMt��+��o�$:rˏ/o.�E˛�u����?���=M�{�;���.:Su�`��1،�~R���&�����`�=NC���hi�R����������Gv7���౸��"�!��T�n��d�R���B�Vf�&�����q}��ŒN��l�H�2K�f�7��MX$-u;}�'D���@��F4S_���Da�,���l�Q���$�>�*�E�Z��o�F�k�P�zR�r4�v,�{K��oa9�=7$v�J4N�󯰽��&`���B#�v-ejo�,[퉥��H#��f�����S=8�98��|䉮�Ye�M9{�����?�8����82B�b��5��%Y����aTJd����:Rt���+_l�2�*�B�&��'���	�i:�1s-瓲�����Q�|��"9a���EW���Ct�-���Ѿ_���ʙd�~exO� UaH�T��t���5Crc��Q���x�r_�8�L��z�B�׆*+74f)F6�P�w�l���W:�,m�Ǥ(Jve!>�uw,#|����^w��$�Y�wP�Y���ss�j����ۣ�;�`�Ok�;�'��G����i���L"wJ� �׫,^!�	{��U�>@��`�� �����g���Dت�'q%B�?C]��!���Z��
Y�����֫�{���/E��kI%1�mV7ΥxP����Г�&�xw��5V ��w�"f4&���,RJ�h��ͺ��������=g�H�/�JJu*SV�����>�y
�6v�r�ll"��1y��]3�9�eR�"U���cjG�,��9�����h�~C�W��W:$�)�e;�����\,hUH?f+	_�a�T�b����`���gQ��WصCH����y�H<<�|�tڛ�d�ް��Aϋ�e�>r3O�cd�G�:�O���I�g�~Lt��^ROȭv�o��W�V��Ѵ%�h��{+�6�f>���y��
��f̜n�e;��h�y9c$?Jp�*�۞|b����z>������;�Ql��iuED��8R��0��.�m\��!ݟ2=7�ޒ�i�O��4]�#���uбН������;�)�y������l��y4ɞ[洏X��i4P�O�yH�*���.�c����@�G5�Wඝ%b拪�[�Ĝ�չ[пw����`,Z����5i6�,V����cʭ6ߛ<D�7��O ������v�F�q�I!��~ǂD�*��cK���iZ5k��e�.o��1��+�iq�?��/���$�cw���	�ف�}�~C�޼x��Pߎ��5��S���B�g�Iw7�yL-r��)/��kaI�L)o˛�w�JYs��F��|́{u3���i�2hLתS.����>�{Y����[���R[�H�Q��������4�j$�-#QՉ669,u\ӠN��:�d�j�a���X��.�"/ ���籌y�?h��M�6��ԣ��u�J|��� Zf�ZSw~V�����sv&�]�p~v)z?TLK!�c(B�MNʙ�Jo�y$���������[r���@ngBK:��W��N��9>��
�q�o�I)*NŌ+ZU���k=�ӥ( �jI&w���xC��gX(ΧD�]�(9R�c� �[`.{��.:g����#�����)���V�{ֹhjT��ʺG�{_"
GӔ֨Z� ��?�q��~�j���x�e�����(2�JU�Af�p�>�����t������AE�������^���!6VjY��1���yc�\Q���Qa�){+;�0J�[G��sOoj�Q�j��N��5رޯX��L�(,�����6rФ���P�$F|}I華"�{)>�Y*�[zi�yd�g��Ҕ������T�7G��S�B��{j��{����<�9W��B�l+<\�+�%���}9���^��[?�u��Y��,�A��"��k�⛣�8 	����э�NEOK6�Y�C<���;�KY���T0��������	��-4��N*j�4I�e�G}p}sB m���׫�+� �iYa���+B��G�c�.% �t�8QS�X��,yg��-������A���-��4���);�����V"�{�!��%������S�^/Q�*�7|�ʮ��0�[32u���rF6���'�֔Ҁ�)7
���w��{#�����sw�I�T��G9��h�Ҷ`�$3n�e��ۢ�Պu9��3���US4�ۨ�+��J��
J.�YW�� `-|��l�ZfP1���wc�	�DLU���+��u�v҂L�p��)GP���7������ �緕���k�ZG�2���f�9���X�d��� �����ݰ����+YK[�ޤf}�����H��2=�X|�i�[')e$V*-<�6MȚ<�Q�'b�|��v(�������b:�S��Ut��QUy+6�%ə\���v��Me�t�:b�����C��$��
��)d�)�����=e�~���m� ]�;��f}Q^��U[�,�ʯ�{ņ����|�/_4~��)	xn����.�`�:M�I8ʵb��Gyg��}��,]�5��/j�5~��Z�@�)��M�sǭ���d�=���b�I����5@�@�;U��*��.ӚC�>��$(#͟;�:�����
;-�'*-�r9�]��=4{�߳  (s�?c��V�o=��I+W�Z�XRz��'�\�Դʘp��� �,+����,s��H	r��m�Y���A,���႐?�7�x*)��7�sMs�$ْ��ZE�%Xs\�.�¨+.-g�YH[7���䫆c��XkHaX�4�i���S9�y����U��1���a�ڻP�ɟ9$X:7��Qׅ����?�ܶ~��:����3��U��\����=�k�я���">�	E�eB�����|��6�>|�l�U�>w L��:sɏX����ܭ����Uf�F�-��*��g��ɝ�}]a�.��JI�'�ud]s򕇸�NJ^����@�U[��Q_�O�D�sq��JX6��8^Q(S20ts="����\M�d�3�����&"�Y���ۗ��|�[�|H�d껙 %���)�&2+b�{�V�/#�?��{�1�K�Ԩ{�Dl�ث=�ʨVS.|�1�[��$�h�$hb��Gҙ@�^:m��1xD�� ���#�ϴ'h�Lcc��AW��R����;��I���7KL4�[�S��D;�f6��Hd%
N+&8yK(@X��t���뫳$�]�;�C�r���G�Y���C����|Lg���:��;c���8��z�郖<��aS����"���NT�kl|H;��ө[@�i���nr�2ST������C�;��ț�d8��ο2�Jn��.�k�VH���P�F��?��[:�r5n��Fc��ǯ�D���a�"1P���&lD�{㦘mZ">;�N�pC83�F极�,�B��\.p�f8�EhG}�yr���)��W׊F�[�=`����N@X��n��dz7V�����Xn��)�K��]����b�s-ȇ���!b#Wi�/���eކk����,���0����T��Ӕbr����-�X������u�H"%Z����`����<
�SoV �y�uY��d�<�/������k��H�)OՋ"Y��=dp/mYxsqe��a�z��@s4}�����-��=�۪�]PR��n��3��<��o�(�8q����H��9AJ��0���^���\d[Y��*�1��}��:�n���g�4o�@6Hwri�'c&�������}5B[�)�O۹�U#�"ᖜ�j��� � ��~��-x�-�;^�i�O��X�����C=f��\��� r�tӢ�M�B@���tN�iJ��}�<����ob��G}+���*��:}��E&���f����Ui:�YC�!��jf�	N5"���!��Z�_�o4 �L�+�{�
y>ʣF�ơN��M��x���*#?1Rd��]��'�P����g�	�#������/����K���ic��,�9P���n�垀��w���-;3��[�ni���;�1��\Ee��,E���H����Y����G�CZǒP�$5�l����i��k�+����c�Ǿ�g(�W�B�7`��l��rv���j��g[(�R(�����(���q&'J��n��&��k�<�4.c�'�!O�0L�l�R'����;��k��y|hI�G�T��`+�������.0��OP��&1*�?%\%s��۬�Q�ߜ���d6 ����ؤyZ��!��pe���%1J9Ӫ�ʮ��K�[v5䍽��hj'YαjJ?�&����&Ŷ���{�+��l%C/[9���Ai��t}D88@�?�,�k�SsMș�K������\{��ިM�ہM��&<�Z�ѷT�4�e���Z��DplM�8O��䳽>L>�2l��Ꝧ*��
c���g�Ȧ0Y�]����ں�
t�m�1B8��*�ՠ�q��Xs&��\,�Z�4�8�v��}�=��JF8f��wj�U�-)��� ~�������E�̜�_*�|�0�v�4���d�ڼ�}S�XNN:�88�?��8[�Y��-J(����!k�J!,�iP�1?1��x�y�&�7�,���hL�5/D���bB�K��g��\'�$i����-$R>�Ϻ�b�C\�����ۃ�u��[�_i�-k	�4�%3$3�ٷrz�q�?1�~�_u���p�� `.���>R�j+u���>_���Q��i����.�G.S$�:Ԭ�\�Dˉ ��?���Oc�������!}z��ʊ��|-���c}��zW���=�K�������e)G!�Tk��-����1���n4T:i��7i�5o��'�_b�c�晔��'��GT��Pw��3��{}j��0���I�gĖ�ܖ�NO�	��w��l�B�㏉τ��官��z_�F��l���dk�6�7d���%�c5ůd�b�����%� �Hka��XO_K��z�����Du+Yp�y�Lm�����W<P�^�SBP���<�N��LWE/�Y,�̰T� .wy��62��y����j�����:z�f&�A���t;��{0f�L�
tW
�&��&r��_���"a�Ug�c�,S�Cfr
I�������D�F�Xx�����/���ea�<�TMF�'RjC�OR�i����G%Q��?��v���OY�
��p�ýg�¬,�|���|oA��6�J�}@m�A�7��K��Ȟ�7���H���d9��ȠD��:~빰j^��R�20�UQ�4���a���9��ߕ��?�L�rDǃ����tQʢ-}�	 Aj��j���Lųw�溷��� ���Z�=q{�P��|�3�%�+jm��#u�H�:	�O ���a���%)~n��\	�w�2��+��W��7!2�I�3�S�!�������g���H�F�=���� �p7[���
�m�}L�wdO�ǲ+�Z9>��G��ʌ���\�e#R ^�HvQ��ɴNi�ý0/��A��Q�u�Fw˘����Xk��H����İo�&u�gXߴ�׈�Z�s$t0�dw���*X��ːp��t����"�ɢ����Z���Ьx�үQ;)��K#�ϵ��>V��Ѝ�]���"�%�H���B�s��QWsT�#,�����r��W�hu=d?#$Y�	�yGA��3y/��X��N� ��2��K!� d(7���#fo�%l�ؑ�)�ĺi���G��x���l����/�u�_p��Z�.�%(e��K�͌��rh�W��3�t�-\*#�-j�·��v�߿���O��]�����Q�-�},��C��ݗ�n(�D����1�:N��h��{�Ő��&2��mRO���gY&�ᱮu�W�<��M�ǚ�͗_�´�*� �5tDMʴ��{����w`�}ӂ�s�P������n)��zЩ p��2�?�uw'�[j�7\�"ؼ�x����,-[/L�.`<�s.�x����@�wX��֢q̱���zK"�a��;��}]���C�+��%nN�=K���z
 <�C��j@t jʂOǄ�o�T9���Y�*L�H� � ���58<Q44���~�NG5�J�Sy��%�h.s�o��pO���F���g�����K�ʶ�Ξǀ[[���4�[̝�χ"=qGxN��%5]���U�@��� �0�$���G�2�&�,K�U}���/�����
��H��z�r��vdl���1�B�������|�:J��-�(T� �6�o�7�	>0կ�D"0�`��ns�$ D>(�{�-���	4�:K� ���4}�U1JJf8:KX�ǡ<�u������I�jYVY�)(k,ˑ,mF.��S�z��*���_��yNV��U)o��t�n�����b�/j��$M��<�Q�	��	}���dw;�qHC��GIǚ�Z�&ZJ�ѝ�ݥ9��!^� ���Ҍ�M�C�VC�5,�a�y������{�V_0��Q���˕f{�P�>o����P��8�p���Y��ʎ�~�K�|�$�nz�D��W�8R����M�(\`TS���R�d݃n�׎�xDҔ(���$��.�0d�LV~��ȓ�U�ӧ�"��S�*��rv��L���J���cW]�����}���v&�/܋�3P���2�w1�r�d}���8�V"����U�srG#F����N�왽��B��7�`Q���۴�8���f�_p��uf C���w��.��~s(0)����X�e.]nw��w��*��d����@�8�/V�%�`܀?�]K������ pp��z��Q�s<��mܾe�h�!����z��|gbk���o�uu�_?Oġ��*��\*pG�BL������ߘ.��LD}T^�X���X�1��� V�+��3��0֎�_k�TC������I=3/rs���&mTcۂ���V?-ϕ`d�b���.�L�̮�c���4d`���[L��%�ʵE���G�ȜZ ��'�]�a�/V�3g��)O�\ep�4��3�L/���d*�Uq�������"p�eP�
:P�z��`	Tp0F��
�D���T7];:�>hӆcS�KU�%��2�Ll�����@yF��ߩ����@�u�G�C{���N0�؄�H c��K��$�I��y�7G³�d�ub!�"��)A�����C�B�x�z:���M7��櫘�.VO>	[��_ե�]ց(ؽXǱ^秠��,A�2?T���8�ב��K�eu�M���zv"S�ױ�\h�ə�@I]��ct$�(A9�a����d/�Nt캟	��� �}BU)*aݬ���1������\�d��k_y!/�㌈�J�"t��"]�Փ�e��?t��M�'%&�������2�z/"{6q��gm�j�1��g4��SجR�@�����-iҁ3���?LG�vE�2ډ�{��h|dض)����j23W�v[�鷎��Ι��g�z:k>�1h��McV4��:��PW�L�n�agpo��>~�Y*ۯKT�����?J�M�Iq$��b����sA����xNCw
�.�� ?{'P��"Ќ��������\�e�l�-k�rѩ�� »
_�%\#x���~\dX�Fs���Oo�_��(�:�F��@&���;��䔮M��S��Ս'FØ���?֒F��I������⒄�����z|�r�t�hf/�p0k\�#χ�<f�V��@E<5�ƒX'F%�-�J�ڗOcgu0I���<����:	NOF�c����HV[�Rf!h�J�
��	/z�] �,o�Z?h|i��e���j�G2E̖��w����w]��3#o�"�l4����Dh�xǇ�A�:.p��b7" �6,w�<� GZ�0\[��u{� �
��X�@�OӪT	�g�B)1g�Q��੪k\��+��{�F�,IB���-�k��X��-���1����~as�*�
�SNw�	��y��JE^�IO���6�������Gb��Sl�'�_����I��s^�G���24T�ԋN����>��8`9w����y��!�Ih�2�ty���J�u"��������Y:�_�{�}����⡤���[�I�A�b� ۄb��qM�����>�6���<��j$|�[q�L�GY��"�J5�#sKڐ@j�	�Y@��F�1$��۝�Je�	MU�ț��(��e�:�r\<.���=�2ja�4�M�_[U�����3��j���;��5�V&���LK%	J_��/�����5�j&�����_�La�mU���1A�\%[:�i)d�J�P�6gll�E��H�6�'=��Lp��#�*�8ۀ��?�h4��F���m@�#�����D��<�0�XCh��0�*���U�L��+s����H�t���s	��z�^�(�'z��L�PD�Q�Dp{W0�h�5"�!�*T��s��,n9^L����%�FZ�4.���N=c�	�g�+ <�u:�6h��5Q�d{�r��h�.��P��s��%H;�}��4{���$�l��C>�ܢ��0�
��Gh?I�,Ww}Ѯ�}�{��Km��v��4� ��@Y��D����B���:� \��`#g?>��I��o��Iৌd\��WUwt]�E�P�p��54���{���e��N����}lZ���?�}����.E~���!q��!L$:������#�=����p�
Q�C})8c���n<}2``mf����w���	*.���]SqzoD�3�"�Pq����֜�~�-ΜD��L�
h�ז�M~�W��v�����e�']�#S���P���J0G��*�S�xs��R��d+c��YJnJ�����G)R��-/l%�R�ܐn!�:�[�����\�;�P�y�3�	�,����{�����k�L�f��sC���T�W�3^ZS��y��_>�,�^>�8�vj��?;�T��.j}�f������=act&sv�  pA�*�1����a�ʙ�;�譧.p�,H��Jaey�EG���.�j�������>�$-�;%cm�_�)Ҍz�� �5qF���/
[���&Q��8�EÔ����k��`�LsFX��Ng�sB$��-�۞��%������%��:bL+Q4��򼠏!_����յ;�|Y�)#��UB����-�{�y�bz�8F1�%��ˈ#]t�L��� �ZJ\MH��� ��ϻ.{��D<~��Z����iS<Z�Ȉ7�AZ�J�W9�2�ޝ���h�@�s�H�E�A����~"h�¯�ZK#z>�9���U��!M��<Y�R�#������)���r�C����E��:�3��L����)�ݦ�kc�r(W�����xj����Vx��n��r���C^�9�ؕ��/���b5,�W��Vv��xɤ;2�*-�gؾ��`?�����ly��	���
ԛ���.��&��_'cT��\}!���q��jS�~i�.`XH#���}3�F<��y2����jʾ��om�_����_���Ӣ���d���}l-n�$1:_Z.'w[�)iZ>��I�[�v���>�+;��:�}йј�������Gw�"p�pRq�*�f�6E�~iB>H�q��$�ph��rY�6ʹ�$�\%�~Lˌ�� V|ȉ���!Z�A@�)k��{��W,�&�f�<�?g�W������ÈD��Th[�kP�_���5�-��T�����y	d:>���8����~28`/����L�%9�-��
���z]��>��xdڑ���9$�s�L^RmM-C��;,�V��=+Zy�Ww���!��&Y����Ҧ"�j-E󚻂7��Wrh������fݴ�b�0��F���UDi�l;j��z��.���@'�Ji\ZC�0�k��>���������S5��{].�� ��t J*���Y��}��^�N�4�����'ȋ�x�\D��#y�+�%���S;0	5q%E��b�_>�,Zem����ɓD�icmyd������
�&�,�7[Ĵ�n	1}"��[���9"������k�b��ݿpK����QEb���t٦����LHݿ��X�%,P�� �7	rm)[��S'�z�9@���<.�o���	x�K����˫N�V�hTw�����$��,}�W�7�;�-L���*��M�)�����zkX��/��+�i=6қU�A�Y���/c��.h=D��9J���)-i
.9Y#��!T���T���G0a7r[կ�Y�����pGK�K�W�5�-���^B*xf����f�yOT�c��0�'��Wqx�I�e�;�<�~n����˨,���m�3�?	����Z��Cw �\8�:�A ��@Rq[��͎8�J�K;?��GA�N�\߷�S��SǍΫ��.o�cl�K_��Q�	p���x�ռ���"�7���(��a![1Wdڌ�S��
��%��3�jMoh�>�s�^ǌ��2Dbٻ�)[L0��y�-�MX}B�i��!���p��o�L��#YB��=���5[��Q1��VnM��r�;==U$�6�4 �@":�/[���M��	��A��H%��w7k��to�Ʉr�Zga5ór���8��#)��������sU�<�<��r�g
�t��l0��64l����d��N��1I[L���tC��I��(6ZmN�ҌG$�\x,���NQc<��%#�_���?�8|���o��'1��������FwYM-����H_��ˑbO��U�>����2U�Jڽ�`��b[K���&e����&��Ldy��@���3V@I�Y*L��AFH�@����vS�q7:�hS��t]���"c��w��r���+"�?J��s����xz[s�C,C|t&~.&��4�!���3��}S�O5٥����*����M�"m��pn����d
����*<���(:mE�Wg]�3>t�`�eT��%�aVZ@�C�97�;����{k������r�{'���Zҕj����w���Nw�V��6�
��>(�PO��*�?���������q?c��"ص���T��Mj'�|����4����V3P��]v�&7�W��Qc�:f�e+ꤽ�J��1�F���p9iȑ/�]�xWS���*�q2IB���2��jɤ���$l��3j[���ꀄ\�pl�B�$��%fı#S�R��Ū� N�//��Al1�3�r�]$�zx'|l�-�s�J��8�=��9���`e�\�<!3�Uݱc�:�r�����*��jRa�4:N�!�FGN�)�$�f��dIdֈV`�#ݷ�l���S����X)I����e@,��g�"=�����z�~nC34�ZQ�&�@)qO�K��7��Zs_���!�
�#R�U볟Z�JB�]g�����0GG��Z</$����� ����\�XR
)d?X�2Q�����f)L��O,�k1�O�Cy���362�j�bo^8ľM�GJ<#'������S�1�g縡�R#��
mw{ĶM�v�)þȽq��Z���:��4����w@Y^=#�(��(� �kkN���D��\KQ>=p�i���t+6�K7`��Y�y{�Y�J�ȏ����5�=������¸�}B���5�g���>�x*i�
IYg�Zޤ񈕿yA��k]]�**���x�^�x/n��a�{_��o�w����xg��;��R0���������[0nG��,�'%�����3�#C�gb�Oj@�|��b���+����u�єE&C!Hm�{�6"wӰe���;����n�~��%2Cɗ(,��d�#e�P��{#�nqD�M���I�evO`���!�5�R��i����B�{�e�i�D�D�U���|�=K$���7������*�b'���t+�[&��g�r"�h��������f�Pq\_C���%������������h��� ��f����2��F�/1w��N��h,�W#����;z����p�97��U���,�czT�0u������ȗ��'�T#��=F�9�c�w�PI3kC^*JtDK��#_p�hG����-NT_�#Ŧ�P�@��EP>��Ǡ�@�,;��K=^,��Ō>L�
s�Hf�F�D����2�u(	v%�����ײPf�ׄ��b���cN/�)���Vʎ��ئ��OQ��p�	�i1R�Cu�Х��d�+{V��Y(��2�u��x�wXu�虍o�������^�<��R
t&����s�6���i0Q��z��e64p��HB��~)YQ�.��ÞE!H^!8o�\G��x�w#��n������'ba\Qq�My씪��V����2�K�d���ѹF����o%����_���x��6W�U��O���[ko�7F��TRߌ�⦀?X��T�ǚ�P]���P2Ny�Mܳ~,�"-�:��^�jdMo����1�r���P�<�e�G�Yԣ�D
n�G�E��V��U�ܒݬ~xr���p�H�0�^'M��F�n���?۷@exr/�iO]3b8M�u?�Bdj�n��ΚV����`/��3�G���5-�ơ��q�<=����b"/ &�����2]�W����jUU_X���Qύ#v��~fJ�I��k�۫���wy65�q�m��~:ݓ�g�b>���hg��=�x8�]�Ig��<���c'�U�ة4	��κ5��?����oT��K�	�	�CBU*�Z{�o9G]{�'�/��ʻ�"���|Y3$?�v�@��E�b$��9�yZ�
�s��d_��Ӆ��qu��-���د1����i��V�G��/��'bs�c���ڒ���#�s?W�Ų�>A@��t�F`R�)6�/�^<p��D��E ��c)/+��7)m���y��'5=�#�)J�s=K��Hh/l�N@��[{0�u�c����h�����F�A'�FCF܇k�7�M���!�D�3Hh��H��%'�n�5�ӗ��4A�9�D�~T*�z�y���>D4yZ�%[=����� �u$g����� �m��;�=�6J�h�*�f/��VF;��~)qun��u�e�K��sc�ٜ�}0��Og��@���R�-;g�G�+`�"��p[8xJ-Md��-;� ��q�ٯ��H�hq�z��V��2��e?N�j&�|U��b�K>��=Yj�>��p����u���4dK�%�M��E� @����G_����!��Q��Kv:�V���
`�i���t��ko��wY���dh�� �k8�0#y՟����B�[��E�
r�k�:ˋ,q��I���/O'N}J����G�.6��n-�x��:L7���q�����=�DY���� �$�E��QJ�y�:�0��^MJ�C.�s���J�=%g�v��/����2́�9������%�v�?'�%DC����"tE�łƛ���J���:(_O�g^��9w�^׏����ħ[��kB��n�&��H��8�s&�����U:��Hw���d�ƪ������̭�b�fc��s�-�է
�Ӄ���J�xl~��R4g:���|M���^��-��a�azZy�H�d�ޛHG'v�W�6�`j���y�w��|RU�&B�Lea��A^mt�#���E�ѱB��@�v����P<m�&ِkѷ�9��x�=v͂ٗ�dʤ(F؅w���MY\�\	�Rm�ٔ�_ű�D�ͅv^�m�$��L�篗���I���2��������!3�z�k���NO�$`c�a<b����욞y�)nn�ޡW��Yo�J�3E��!{��7�K�$�,�w��83c2�k�O�J��KW}Qq�s�2/�]�1�Θ�%Pϙw-&�G�I	;��Թ����hI��zWg�/+Fa��<�Ѓ��X"o�,�DQ:��E�!9|�!�=�t� �"f�^ق̒7���1#���`��F���Ā���\����Y�i4��"u����[A��m�D5��'�yĬ���'mD�<j����#D�˚A�e�z���B�!��8&bE�D�F��Pe79�_���Z�*�(�a&li���D@�ǹ���N��n�h�Q �>��tS���z�u�T:Y\��]'��YQI�����
G��!D���n����X��������%���i=k�2h�Y[����}��1>0:͡��dՖ³����������0M,���?��5	��g�$b؅��m?g\�|d��0�%/3��w|Jv�.P�ܭE r��tQ����X�ɚ]����	���������` 3��fJъx���T���:��T��n�!�2�٬��cɠ�vA�*�Q<*L��uV���x�qY�h(�FhlW}�6$R��f������8`♤k/X=���Ԫ�`��;a�O&��Jl��JB�	��K���Ӵ�f+ϯD�2��G���cԌ����|f��~M�9h��VE�����[w�Q=�yd{� QתFڥ��;�1�q�����p��]�ઉ��X����ᨅ߿�2n\a@�~�%�9�� ���eJ��@�Il|i���~D�!U��	����H�a��i�B)���@5�>��4�я�q��	��_,�w\��6���ЫHo��>ہ@��݉e�21Q����6Z�-ױ��&���z�<�
��-q�V$ʌ�1��(��)�`���ǽ9@#��2~�dNsLC���m���J�W,��������Tw���bP�Iqx�1�d�{��Bƽ?��Lڸs͒���IO�
����+D:��O��Y�á;<z;��1��ժ�>�p�m�x>zN�x��x�{�[����?{:y7�pF��)����L~�)}���c(1�>1`l�!���<�'�K�nS&�K]���fP��G�m]����;3g9*ML{����2�J�y^
(ID�#�1�մ7�
�K�N�f<�(�\!jO�پ��#C��b%�Osh���E����"[rJ����CplK�|�&�":j�·�в:9�����1s(
N�2��tf.(��r@�K��L]�#V_	���wN	���Z�����pX�m9
1\��]a	bw�+Y	'��3��?/M��NN���"h���!E����zqj�ߡ,�� �p�u,��6�3J
̝���x�Vi2�����y�d�lڕ�f�	U�V������p�`��,�gH'B�
�5����X了4��G�e�x�*ĲVi��7}\��ϲ7�4����r!p8���L��^��f�0�a�:�mw�s���3�+..t|��H!V8�N�hD�X@v��_k�(!�ts��l�D���R���R��ZiOr�_\��1WՈ,���!���O=�� ��Nr�7�1ϔ�M�7sJ�$�%`7%��΍��m[���oi(f�S�.8�g"6�Mv�Q��̆����[<�����vޏ3��S!m]ҧ�٣=>�n�و�	���A�S�&��Kj�\|��v���mOCn�%��
��s����S[��b"��Ĩ 4�B�!:3Dz����iy~e^�x������j���I&޵��"+noz/��oZ�1�;��M�,hT��{����0;��>�	9��L���W�0{6��&�g�n����r��-��l��#㴂������g)��\�֨�D� u17p�������d*X, ���61�H·1��}9�M\7��,��.�O�h�i����/��F��/�z@�?����֗�|����D���Nt�O&:I���ow�9�w�&�z��� ��f�lv0k �� d���$ �����
���c��='H�E���L�LI�(
�3��c��h����{:L֢�*=o��n�M���Z��6��캂2��Wx��NB����X���`]Y�P��P5�J���j�M`x��5�;��q;��jX9��P.|�C
�O����I0#S�^옸���M�6�V��䵯�C?��Rk�$�>"��=%Z����}59_}T>w�r(���4�DE0PIE�y��x�M;��������a0�Z��c�'�*d<�%�}�� J�kpF��R$�n�٫�.�a�,�^�d�k��d��CS�W"٣l�'c��Ȇ�������:Tpw��6�%d�����9�X���{�6�oL�'�����~���ͧH/��m^�"N�)���.�vorE����q5pZg�c
�Dy}AUo*M��x��D3D�眪Y��u�jVN��9,:�ȣnȱ����M�	m��඲)�ܳ�R!>:m3�>$K[{_o�+���!J���j�������*2xMu�چ�w��Ge��#H?.�<a���t!���4��%�}�d�۵~3�je�)^�7`Xy��b���_�if�8�s�L<�b� zA�n��S4��0����Z�^sH�D�����w���ej�bv�`4��6h�"����}�=������Q�T�q���O�*e�%N��u�)3���؜�5��$�d�{�j�0�^51D��t���su7��,�~��t��ʣ3�s<8t��^�#��%�d�_4-_y��8�Ba+}�r�k��Y��оe ^��/�|����LA��x��x&r�Xv_�]|˸�4 d<���.yϡ����/Qi�%�z@3e5m�Ԉ����ʳ�sXPd榫�>:�:�W���M1��{Z��MF��O��}YG���:�7'{��h�*r�b4O��sͱX�Hۢ�Q��+���D���B\���6K6[ܱﾔ�����զx5�/�-����cО��ڡ�"�0��j�` s���e��fN%(1q������ƍ�7�V��`�f<�.9�ZU��z�q9\�h�����W{�._�Wz-`���ѓ6>^f��لd�y��K\5%f\�<D�t�Ԗ����A�*�^ߩ�����;d���/Q.Q
�]n���nke��fПj�[,o���O�x/��*f/��_��1����G%�p�?Ob�د#3j�;M���}ʰ�����ի���cu) �3��-m��S�f�A~�*���éj8�f�U��� {��(*��x��5���[l��3�S����� 7��b?�s,I�`2�`�m�"yF�
��`������xo��*�wj�4�Ve׃�e�볫u#��I�d�&U�U�����v��Y�{�Eߩ��}�te����z޳MJSg�n-��6��<r���kw��!J\���]�ջ`��YV�z�s7�AYV��kH������I����~Vb��yz�3���q�{���z*��_�T�Ӹ��޴���c��xv����6���y����zl�2�r�(��4�=zf��g�����<|������^^��@J�΢^����]*��'��+�`~��;�m[��~Z��)�q����QC�z�?�[L���qD)��d>�}���[��Ǒ�tK��"�v��B�����p�o�f`��ɦwz	4��2ȵ�A�u�����so��J�aJճ�+
t}�$��և��#͡j���'k�b��7:���I.��&��UK������}x����E�-P���w�fOǉ��C� 8H͝i ~=���'J�=��_M�v���C��>�:{/��W�������~siyC?����I���|�c�ŉ�h�a�lr4��d�x�����l���L^YF�&��_2WsEl������]�8S�Y8���f��_6</S�Z��|���/Wk��1�n���%�����_�n�h���ń���h^�\v>bq��C"W�;����Ux�9��>�<�/���w�|�*���$#ΒR�w ��M/|0=t��i�Q�C�� B���q���V�i䐸$�u�t��8�WqJ�sv��u�P2���Uj_..3ܚ!�%j��C�H1����>tA�s-�}fq7����	�Mc
�/io!aca��&#ӧ��_(
�Mp��.��&,c��AA�%���;F��M
��ߔ�K�/R�x� ��o�_Q�J>�m��n���������g���N�h�ܱ�{K+� �t�n!�[%�10���$,���cd��Y�� �x(j�;�:��`��)�?����	���Jpd{����*��������e):��@5��
�\�c�����NmC7u�8���P�oh�ܵ��ؑ�l�q�ff��@��Sk������U6�(��-�T93W�����2]��<���&��XZA�'lPN{3������^�� �^��02Ow�X����bfT�?YumQ��!8dD�F��PF���N]��7��E��B�����r�H���{x��Ɓ�"����S���b?�e3��u=5�)+	F{�\H�o�H�-�h=�m�r�|����b�>�����z$ X��(���"Z��:S꽰�#y��⮢�A��vP�l]>�Z�1p�����?+��v]�r�j{�mS��D��ʍ�&��L���PHc��6>��R���1�~'�hGDQL���p�L�zC�퓧J��3��WJҤ�����	Ԉ��,����.�	�ZkT�o:��|R��\��
D� \8��i��T����`���Цp�FfQZέ�>L*Iqy0<�`2\��=u�T�W����5A�H�hA�tmXkȱ��ָY�5Y�̀�v���GR|�n��+@�iʰJk}�!ķ�)^~�z��1��b&�h!�,�Z���-���X\Q͋�Q�R����R.x�M�@������ޚ{�QQ���)���Tl���O�aYH6�T�a��X�e���1F�f����|c"�&7�RS(	����$@i_}���B.d��1�続Gn}_�1�.0o�[{Zm�β.�a�NO��f��o��˹�&���
�op_ ����4��9���!ʆ���J3<\\�L��W���]���:�$��P�[�f�/A��F<��kE�Vǚ���\�-.ð�"o���bЕ�V��%�Xk/�_�����>��F\0y��hG(��2DWlp*�Yk/��R��]���A�TmL�@ԙ�@��0�7ҝ�2)O淝vr�_����q�M����=�Q��B� ���x�FBO�ѡ��i�������)4r�`,|��u��������UH�Z(�-���4 ���|c�)"���{�WS�P��:������W�lC��=�,��g	����e^��Bz�tR�^f܁QR����c�+�e)��	3��ñ<�I��(�b.l�:�)�&~i�륔�AaN�H��4[�y�*���݈�7��F���k�A�����w�U�����씱��'9����K���� ��	O	u�Ħ� Q�eH,'��kh.��)���4�?E��]����&g�R;̝r]%8|j�B\}��:Z�;���"�Q$v��1��,��ο s+N�|��b ݶ�&��-���-�m��6!|�\hӻ��2��㶂����f�fс&;^���F�δ��m3��[���5�C���XM-�ѳ��R�^���a��}��h��9�uL'ON?��H�a]Ȩ�b}�J+DxM��������i>����{9�b^�.���5-e�� �AM���u���(��$����FB����]Ŕ���1�\"8�6��݀c6i򤥾����>D+J����$Tt?n=�#��vr�N=#�y/����D0ir`��)h�	a%]T�C�9�oPt�b�,�F���A> u$��_�6�$57c�~'^H	z��e}�ETQ�"F��cbE x���3my���Ȑ� ��c��(�X�@��dR�m4��d���BX��t�z������J]��@���С�}t��A�K�Թ�*������)�f�̇��ד�,M�u,&�*S�!��:�t�R��4�8}P$���ŏݪ�F��I(��J�,}��]��F.�(��{�bm�2��
�f�n������F�t+7��a�mNcÏ@���5jZ�L�w@\���ldu�����o��(	]C�A�n�X?�w��׵C~( ��[`��ћ��y��n�.��%ޟ�&DEG�EZ|h[�� g�.��Ϸᔗe��_L��Z}�V�u�ic��9��Oۛ4�������di/o�����ů��_�t8C��	��F��Q�g-����ͳ�д�WG
gk��/�9w?�r+-DΉ��%�9p��w��8e$<���@��Z�k��K���O��nΖ��GU������� 7���P��V7�Ƴ�0������@1�{�P�B��X�U����/�����:&���gb�#F�B��t��mq�5S�\_̤��v�R��l��֠�ܶI��N��}����()�|{�,����l�Scİ�F�i�{Mh䨊�/ڦ_���b�,��*�Wy�	W%�Y��M��'�u��<��]�QhU͂���^��A$4�L
wm9b�|�;]����R��r�Z|S�����ܶ�pa�=*|�-�4xBiz�J��(;f�L���4u�?&�G�UЃ=��h����c�8h9Ŀ�0^����pףc��6��Z����-~�ZE'B�!s~��u'z���/3������a~D(m���K�������[&��K�o��������B}`�����r�w�ѧG��Qy�������$.~BL���h�)g�g�$�u]b�SN[A޹ O��&ءV�j��שbju�f#�0��*�V�^=�ʰ�^�L��Z�^��&�l<BY:ॳ�7�ǩ*���iq���>g�X��`!��+�M�n�`�ZD�̀��!�c#�b��$﷭#���6��Q[���ٯ
4L�7E}d��b�W��Ư�yG]4Дv�����y\D�����uM��]̳:�P
q�T���3 W�?{=*�%۞��͓=8��j�A�m�)>(�+ӏ?m�\��+������sn%F���)��ԙ�Z�#X�IG9Iv��x��ė��S2�3~�'���7^��Z��x��Y����g�ĥ�v�9��?;��s��2WҠG��ksU��&��ùխЋLXÀ�Z
뚕����E�92L;娙+#x�x����MҊ�ā��D�c�	_Ft�[!,e���W��|Cj������_m����\�`�x�" �r��0a���J���=`��;4���5�t��+Y�VL�BVI�r��bJ�3f}v�5���Ѣ*I}�tݐ��a���Ls�b<@b�S����qE7���7�]��*��F�](b�0d@�!�.����`���^�����{�t]0#�u��A��z@�����W�)Z��I�~T-\���<�_�;QqA��2n9� �o��s����C�I�;Ҡ��-2�X�f�9��=Ɩ�1!zi�m{T�Si�)N'>p83A����zl댤?U���E?����ӌ#p��N}�%����t����������(��>���g����u����K��h2X�w�p�K�Y t�2��#O7Čq�6t���]��10-���)h�/�ͣ��7�U��x1	&�z6��z$h'�������I�DiLjW,� sE7�u�0,� >s1��)Z@C���AԹ�WMJ*��R_{���"%$�s�ו��8�oM��ʚ��ׄ����,�|��G������;Y�J�R�L4�r�!�a9B+��r`bH?�l�j��醅���d����"�x{Ѻ����w;��?#�HX�����>��K���I�.z`߁쩰���m*x�@8�6�= ؚE�b��{������o|iR��6�wUh��W�El�.��fކ)�*�ĊC���v2�hV���,,H�ͯ��5�s�L���st#�����"����"��s�i���U��>����(��{p�=]���B$-w�'I����͑ \�
�	0�!T�Va\ey�_k9�O;�P����t��h���L��8Ā��Gk�o�~(��]�HN��ϐ��N�d���FI���5+1t�xu)�*��.o��C5Z")�mg
j�U�*�8� Ɍ���H���J6ko$��G�@΢�PQ�v��W5�B�k��8�� LI�޹�kh���u\�ΗU_(ּLs#c�}+x�T�q.3�,�2R�2��@t$)=�}��Tő�/X���l����T�;�d}y�	���8�(�`��}�Zw���ψ�?<ґ��2O��U�Y�@�T�a��H��k	ĸ\y*�s��4Y��H��.�a������J_۸�$��HJ{ή]`\=t�=؜�Uu�)7�v2�e�N�.y��8A�q0J�e�(f[�F
6~��K�a��d9���<��x���+\��MG�%��}΃���/q������V^�	��U-���:��*��>4�������d�5��Բ(�/X�xU/�zѕ)�j/��@];\3\��=�S}j-��1��ԋ�m�D�OS?F)���D\ҳ��A>�f�\�ƍt}>,^�>�Ͻ���$b1q$O9]���ΈO��=)";qXpn������տ�;rA�Ӣޒ}D�Ƃ�V���Zӡ�k�W|�hY�+l��#��:�=x�X��g���ܠfLim]�����,�\�����F�K�<17 |�?��3nN�;A�y�`���9�J�{mv9��ծX�Q��a4��Yn,��\}������U�Y�sƢ��5"_[>�<k����i+9A+��>1�;�����[Q$b���T�IĊ��=�un�C�"��q���8��]���s�.w���ER����Dڅ�y���`��C�G`��̇����ݤUE��pQ��=#�^E��ַ�dW
��a�免�J7�8CP�2�?��������">.��!��%��aF� "� ���(���8���r�)�-X�w��V]��m����9����N5�顼�EPk];��@�7|//AYo }���T�����y�t��g�m��}���a'Ų��h��-1�b�"(.�V��&E|6��Q�jHF^�!��ա˺U��ۥ��I�H�y|�0fh8�/��u�&k���T��|�]oh���a�g�.�5�D6���=�wD�rB.��Ok��dgwi]k
��W���⯤z\Oҝ���N�U�4��ܼڡ%���vMAҜ��.�uF��csX� �TF&%&R�?��ǒ�Qi��FI�t�KТ�Q�ϧ���*�o�xU���ߵ�*��-�X�'e��/q�u�EĠ�a|��XB[c_o��D�Y�O%c[�SJ>?W��������������h��Y���W�H�BN���.�F}�R�3�2_�4�7~�1�,l����gTm�OĪ�/j��<�x����Q`p��P�h�gu�,�q�^P�빬������i�R�Tmy_
Hn��[ɻk�@M�m�t��Y��ά8�F%}!�+ޚ��z�Y.�x�@b��wrD���M�,�f�Ϛ~�Ɇ����]����thz�mutM�թY��јx�7'��k���u�=pj8��z�����+Kn����,`4�π:P��70�����=��ؚ#�c�_�$���}:�F@��鯇����g)|���G]����Z�cb]v�j�J��"�CpԚ�f��W��S�ܙ�Ǹ�C�=�Gqa��N��I���2�5�_)��;EB��/$V�FDv�n��
��f�?h��C��=`��j�Rms�0��C,!C�7��*�iV�����GS���w�2���M(.�l����1���&l�Єhtv�>������EHPc��p8��u�����ұ;#���Z�A�Ŝ�_.TtR~&ɗC�Ccg�� �lO�2�lG�X���;�
έN���e��<��^5�w�(&Z�V}����sT�ǩG�f���wy����'m����Sl��"$ĭ����Q֯�H�DU�J��ٟ�؈�\��<n�:�沘���I605��\���Xdc'��Q�(a]��!�x���32~��Q��1��hA�"W�"ox��PpJ$������~���ݽX�~��D�Hs&�x�H,�Kna����tj��������x>�N#1���pS�c�;_q>�'�.Å�P|�|('�I{�|�={;%0\џ�W��PEre�`O�ե�H1�$a�wO�������¼�Z/���S =F�<���Q2�|S�`�oH'9�n�2�bl��qU]:�ov��!�U�돎�h֪�N,����l�W2:�����A7�<[�	x��tr(�P��A�{�	`Y��)��Ц7��àw�YX]����C���&δ�w�[ ��AD�I�5�tL����1��\��\��A�I��;A��Y��j��QKǻJ��&mH���~��"��ķ6�O�_��`����o�:C銣,Z���m��T�>���˜�t*��2$�d�G˹��H5�]�:l��:*��}T���|�lc������"�C�S���׵�lԐ4�{���"�`��d�/��&�`KBlݩ�����r!`���������"�~S]>�;
�����S�{K�7B�U���k�Z���^+t��〛S����Bp�=8�DO�_�z �UA썕�פ.�7p�@z�������(�條Pw$i�F��
;E�Z��չ?��|_���H��8�2B�l������()n1l>�ַ^E�kU\���z�#�����j�&�g���WKwA�k��?vh]Bn�^�Թ�H�>[��e4���wiѯA�Ň(��79�����2L����6�<0D&�i���ɑ4�����Pp��:h鬽X�J��6:���WBfP@�V�0�&ľ G���L�~�BG�Ax���Z}���X���ص  ����ڥû����������$^�9L�_9pX(���1)�0���(�&(�7,e�G����S^�t�*8F&�KߓւҝL�?���El~��+�?���E8zAYl���@���S �i�4�s��>ڸ�n ӍB�K�f�oa2���֮�+��M�q��Ԫ��^ɳ���8���jl�����V�YM����H�g<�jJ���*H��L"̞Cl�&�w|�duTf��i�#��ß�e�s��}\G�l�+�N�/G��4��>���~�-�=9x_����@x!��5ܿ�<�m��g��)�sgkg�i��u�}�0�(�����;Yh��Pj�3����I�1IT�d��k�^p1��C'<��;4oe��a�b�D�E��!�wah �A�O�R��	���-T�@}�Dv
E��F�`��.,O������^�S�>^����� �
`�i�䜗n:-b�x&X��^$,�W��W�CN�+�ݤMSÏ\ �w��q���y	��Q��x3��x��&DP�w���JU����_�s͋x�3=��C8)]JOZ5o��I֡�s� H(�P��lO�pL�D����I3�=v��j�7�K'��2��a�(h��9o�P)햣f�l���%~w��0;E�2�/����4ϑפ�
����#�h.�< n){�Q_��<0�S����H��\�չ�KU)J���A{�<D�g\)�6����ssՏ��\|/�6�ث�WP�?,���S��*���Ք��0��t����I0�	�8����~��ěՇ�lN�]��Q���ۚS��6�Wo�V���O!1]^�X����qsוb�6���c������2�Հ
᪜��|�dΪ"�?YLN*,���?�j�j����LK��p�=?�Q�� <��O��ԛzG�}�2����~�1�)Uf�U� ��1�� ������=ƥ���2��TC3��q�Pօ�E�>��;Tl5�u���um�fi}������HN��4�تU
�{
�$G�T�rkm
�>���*Pf���l�|�/��J���~���'�)vhW����Ø��в�9Czc����;R��.�Z�r���fVs5�u{d�����00��0y*��(ٚ<Q�p,,a��	pY8W��4ޥ�>h�ta�m�	jњqP�7T��n6�U�ˀ)�&�
���5ʒ\��Ά�v�VZ��	��S�E}�?e�JNbp�Y�ș���ߍ 8"�����g �5��4�&-2%W�U����sc_��>]�z㏷[��O1`�R�|ɪ��P%->�o����V��`�ce�p�Ov�k���[�Y��Ђ�&!�;�M�5*��֗���b�u1/�b��޶9	�3������	�4X�f��	�Y�����k��`���cP��z�[�ՐΙ:[��,}�~�XǐJd+����u|�`%@����À�Ƈ��c�u+b�~P�����v�'�W0�IG�t8����vٳ�4f�ѷ�K��|s^L��f�h�øn�����(����$�+�k���E��3|�q�,CP�)n=�=�����.���A�������㡳AR\�6�Ha�|��]-�
�E?J�U	��X�G�e�?&c��{)x��a��\��\!������D�2nTgY�����>���x�_���7OU�RӀ�+�����~�b����O�Ynᕝ/�j����0^*�,�V�b"}�"9QG�)��B��
�@�'���d,�Y�M�Q�QB7/�{e��%�L�,�y�3�E���O�xuM�<���jK��d�I$v�6 [�$� ���/)����~rTд�a+�}��F����;/�
�	�V\� ����X3�>��Pv���_��g��p�5�Ly�)�0������	1�}ߔ�lEp����8�.����Y
9�av�ʁ��g^����_T�>���ؕ�_9�
*��
�LN�f�G��;�+�"�菰p�*��b��M&'i�J���쾴�6�u�|�|�R�V�����%`=�a(�)���'���%��}>��r�E �����F�Uԛ�zd��eN��^_$�M^���� ���gQ�a���UC�8��~���j4j�8P�56m�@��.��[�#��VɊ�#e�h������aJ�+����8��{vB�l(����Nrf�(�|���6�����`���l�{�K���䟓GM!�G;nl��8��dQ/Z�`Q�jLM��Yͦ��ug�Ho�	R¥T�}�>red����b_�����]�����F̗�jjW0����ef�,��
 NP�P�&�.W�_ ��Cu��Q�w<)	� ��Q�L^C�I���!ԕ��1�9��Us�I���?��dL$iߍY�,�7�F���{݊�\>�o�p��`H��g��c(gC�E/��k�J"���#�s��a7�늣�2{&�	"v���V�vtGN%�$I�Lj\~Ĺ�~�d�p�%`���|��b�T,��0Bkw֪ؾ�K>�����͇�!�c̟-P�l� �<�Uv�$�Vj�,:K	��I&�p-$c
[����}	�ƉHh��FiO9Z��%*"1��ި��6���i%@8�a1�!�!��v�$�x7�͌��Wt��_�U�$\-�jU�K�5V��p8�/'Kˆ�(�=��z˘�aC+�"�pK~�]-�i�a�?z�e�y�_�K	`��깺�����҅.>a��P��RKd]�1&)���Hwh0j�N��*/z0�@�D{h�9����2'7Y):��'�w�S(��&����#(�����j��]1�I�F�U1<�Fj�j��ux��KQ�������1�Eڴ�R�̅�Yѐ6q��:�����LJ�D(�ky��kB%�z�|ʄS����Q]8�=�Ꟙm5V4�\U�͡M�P�S[uy��$��i�|���{^7Q����cξ��t7d9�bc�"簇���������F@�B�Hǰ>�"� ��5��\d?��jA�n�����{]��l�m~��4gB��kn~cc��y� ��W�v}����L$���*����<�ۥN� �O(4�Gm�D�}��V�-�Br���7^�5��ULa?��]}�ۦ��팎��C,>j�ڧ2� v�a�0N9�r8`���%�����"U+(�df*ԾJRk7�q�	�c���C�U?�G�!,~�K�n�uj�Ȥ�U	\Y�j3mW[�d�3$@���ii'�`�ߟ�����c��B��� P
i�%�{S>m��=��M�5⣒Y�Q���ԀWOW�+^���W_7�T��m����"�������ŝ��#�X��ഔWcN7���V�q����!kW$C�b~��U`e���h� �O�D2&9��+�㟓4�m����UaM�	!~ϟ7�f��6n�dr�}T���s��m�/b�3���1+)9fy&�o�M�nr�6���0Q�ˢ����4�Fa�t��hKXD���"���=�B���4�/om�H�Mb#{T���kB����Rfc�� \F��~���]�T�_.���_->�6�H�g�;TV�5Bݩ���)�˴9�6��3�V ׻��%Y笮nM�q�B�U}j�x�(���ԧ�K�nl��HK�� ��d�e�4W&����� �\��w��N���8ֺ6�$�NM�??%�q�Ā�"���ݩ�m��&O2�^�1�!�����5��� ����7���zdH�4qe�������qxf7�|u�E6V��KϑEk�Τ�yJ,	�uǶPv�t��� �Q=\��}�3D�n�j����]s�|���Q9�����9�8�!�D$�=Ld��	W|�=Y኎��\��6�J���`���T� ��6���7+b��iwy�N��2�H�P6.*h��\2K���|�#B��Bֈ��k-�X]�(�:�	����	��Q%�A�jL��*]��W��$
?��1 �<�E`%���r�]���^ �����]�o�>�@g�6�F�����|VT�Sכ�",���"�rvG0�P���=R�w���-�t��֋Ɓ�3v�a p�������'O*�ac��4e�w��dh	>;�����&���`/��QZNנ��OA��susF�fȃf�W�LG$��ٮ��^0��+�{��Z6���+�
������y�q�Lh��\��,� �p�Ac6�EvԄ3nL��l �9̌'po"I����Տ����~�Lp��N����r�5������U��圌+�-2&z�V�OߗU�Uf�O�g#Q�2��~���u�������qS6eQ,֐ZC[��Ѝ���ub��H*簋g�Ws����@։#b�Eia���I��",����Ě�	��� ���*��~��ڏ��I�گ�PT��N0�n8\xu<�(-�+���xh˯��`�� =��F�C�����+���@!����t'	<�M�<oX��)<y�<N�����%ІՊ�hR��^�w8;��_�h�&�l��ES�
�b���5/C��+x�p�E��k�����퐒��U"���'
��á7�p/6��u��SAk�Ar�/���*q#b!*�%7%ّa|K��s�k�v��IN=��#N�-�T"�p��h�x��\I<�,%_ ���Lq�S���U<C�����a�*�~���?�n_��ۻ­�X�o��n/�T�9������j>���ݒ�+����Aϳ���-d�tµ�0_�����lj*&Dp$EM�,�dcN�0I�A0��Z��Ǒ���]���,���	B���굣�!)����Y?n˴^9�J�������_j����������i��Ce<;5H����QU|��wlQ�h���{g��'��V4d�WM�ʉL�_e��o������P��r�Yv��;�ȷ��wz����'�+�Y��`�쨴���+��l������1�-P�-��8��o@t�X�i[���Ӑ%J�5�G1��g�b��[��6�½d����#ZDǞ��ϫ M��sF�G�'j9uʦ��$��`]�<�<�
���S���R��JB������q�qI�n�`�-�.�X�.�����y�HB�t�%~Q�V醫�F�1����3		B8�d ���f�NË#�ʐ�~ؐP����k�sg8�+���������v�d9-�X�p�yz;��H��e��L�k�5KlyJ��O��k�y�4|��b�`�v�π�"�c�?���+�Ό�{�~4Wb�A1��KC�Z>��� �+Uj����wK��'�=�c����yQU|��?�:��7.E�e�{ӅԚ��.�]���^��{��ǟk�*ib�:��l�ݾ�T*3m旧4R����3��I�� �T
�x�4����!)8Vh�	IQ5��(�Ʋ/���'�4����cƉ]b3Y񥱰2� ���(Z2���)f2P0�s]7���-b`�n�����z�o�K QcO�v�HI�k�Rėj�2rN=�Tq����B���J����ƚ�isR����ܣ4�?I���!%W�P���Y~̨��R���@�?[%��}�Ă6��,x�pH�/�G%�5��'��Y�Q\&?�j8x"�z�'�$�p����$|_��wFϸ=<��XN�'J�����\l����3�\�%<U��Sl�26��L}�p;x��(}6KP0ؿ�����-�y�G;a���FQ�Xz {���ǰ����I��G�Z9�b>>E����f���mxy�7��Ja���K��������D\���O�n����g�����?R������AEQB�&�wDG�W�ݻ�+_��y�k��&DB�[i�l�TH�`iSb$H�/띭R�]Vs�i��F�l��ҍ˶���=`EM�V
��Ǫ���T�2��tM?\Ǡ6�S�<8����4���a���<��Em���s���\��v�W~$�{�
i�,۝��Z�oQ�ȡ�暈���7� ��~����.#ݛ^��_���Q��^�S�I�#�k��S$ا����(�����rd����ɂ�K+e����0���L7���Ҡ�mÿ}�'s��lj��iz�鉥��[6����9�v��;� �ո)vg�OݷB	�	a�d�)��j�뗈���#��u �=�4Y<b"�%��_#���l�y��~|�Y`��H��������*~�D����T� ^v=�X�ch��X}}d2N-c�|T����핝�>K�l���wb+]dmXy9�Qu踰Xٶ�X�G�5T�H1�,�a�~޴aB�8��JZ�A�:G_�)�ή�8a�/��1)x��s��g���U�s�t:�^	�Ge��Gq?.�M�\k�uW{S�	�E%��A�dZ��[��J����86+���~p=��GED+��=I~�TN��G[�`��+��3$:A�nV�1/�1r�&F?N�"��:�ip��ҵy���������S���[�p,@���}闱,	~sI>X��O����jVeg,+ޝm���� v�xW��77|�:q.0r5$��n�:Uj��/@������V�� �I�a"	�SuX4���_�����J~���������Y�\�:-23�s�Z΂%mo��]o^}��u)�W[t{���kKAÈ���-�%�I�a�X���P}���q;���eEivw83�,�߁M���q*��J��s���Cw���������]�~���whK"��J����ܻ`�\Y���u�}X�� ��4!|#�.5� )j�1����PA�S��׭յ�_ܸL=�W 1Էl�e�\��4[��?Q.OU)�|6ՠ�̐=k�C��?���Gh�?Э�m��+~�}����	g~K\�d9��+�+����ʜ�~�zc� =�\
ûF�{^<,I,5Tx��݄c
k,e�fΦ!&e��QmMT�q���i������kx�qY1|�&*G�?�	���!��z�V���}�-�ZX����U��#�����q7�J�4�@C�Qtp+��E�r@��7y����us�l<�!�˰i>��|ND=�8܏���y��X*�,m*���Q�d����� ���+|0��l�|p �?h����aE������pHW��W����診�e]Gl:eb�%o�q6K=3F�,����OH3&�**`��#��:(i;e]G[�JP�$im��N�ow,rr�t���Q����^<�g��󘇶���z���Ρ�u_6,E󉤉g؈&M�ݖ��1����9�(mى�Anl�h!�u����4��)�F�W�KN ���oi~�0+����W6z����CR6��x
D��^ޣF7�sK���(U.�ˈ8������F�ZU�@�<+��x�d��ed�ǌ���jJV�2��Df�ê;ܪ{��y��m��&�Rh�bդ/���v@�Xe,nj�p��ʨ�F���Rv?��0�`$>�~�Utt���V�7���(����ˡ�[1�ƍ�0)R�.%��Y��S�4�]p쭥a6[5�=��1���^�
@�0x�98�����g��=�,�i�m0��D.�����Zw��X%/|�dP��R%��H��v�6�e��s��2k�x�����J�L)���M��Ӟո���1����hՃw�H�uvbS(#�Flċ� ���	�,�m,��!��ԞV�>���n�pkH�X_P�0~v�q�b<��CV�ve���K\VDܤuc_�3	�k�.vQ�<��މ
,uH���@�Z���z�b�Y����>��d��O[��W�E([)������H���-|u���Ϳə-���Z����B@L���ՙXap�*|e^�r)$&�����Πb�/��^P���En��N|VIޤ�����L�i~�0�.0w|ꀤ�qhkඳ(�ȥ���h�Y.%5+���>�s�B������]x��û�D�}�/B�3Uh��u!sI�t}
��}	\@;o	�i�5��wPs�J�b(�n��mPav4�|Q:33�̡yw�P�
E�i����B��2OWW�Q���J;/̅(X`��*C �����2�gR�	�6S ������Ca�����bI�+v_��nV�{̽�#�f1�P-!��qz��l霌�o}ø�����������"��\���BL��B��3�}�Y�D	R�8�x�����Y_\��J%Msȝu���pձ��6��� s���%S��d�C��c�V'��Lw����F!�2c0�~k��<?�&Q�cn�XrZ����_������@?+��5�A�\'�M���$QG��w#	N@#�Nu��A\���"�\��D��-�#z�iK����S�9Ā�%z�F;�����a3�4ai3��'ϊxJ��)��y�u�	�K��1��S�޼���)�(o�Y���>�U:�B<� �t�J�/_T�E�L?~���{���$Uu��:zlh ����F�ܤ���ɣ�����?d�W7$�o�����b�
X+��A=�bW�)R��\^t��"p�����-,X]K#]m7S��{�?�P��x[�Ӫq��'[m��NbxA�9$�P-��3�:�A�N��˂呃�
��ad���AS�� ���)u�{��A�������u8�G��-�]��!����wLB���u��߼e�E/4�`H>�u7�\vn�]Df����CA�;l}!���N9/nP���9�'L�aM�ӫ�;�!���r�VK?�:F̣���ިv�=L<�^_Tu6��Jԫ{ ��F��u�¤G��{J�I��Rn�U�$'e �aժ���G8y�n�P7�$��I�0��X�h�W����lB�~��Nլ�i��@3�}��(}��T,�D�E�"k<�	.4�wq&<�Ρ�ˆ�T= ��y��!:��?K:=��=�n�������^�9���c��*}�y�}��WM���@z]{&�n[y�nkϪ��0��vm�ҭi��A�3"Vv	������$ƾG	�����qD<I�^���m;�*�l���Q��q�cq�q�A�vo��q��"zP�7I7G�����o�� ] 'Ƅ<:���ؙ�Nr�Z�Γ�V �;�H%���j'��*w^�B��{���+B�d{@�;?��[ee�w�2`�����B� AЪH;W��#���Y��;w�qB�m���hO	.U�H�y}�j�[&�����Ž��/�.J�# �_ޘ�(-���<gD�l��fXa,��3�N~O�FG�d�-֠������.0�}#�yX< 74�ƣN�F�<~�.�o�fX�tz�_# %a�?�������YKi���}��Ն'��EL���Px8�y�љ��[3�S!>d���;T�W�!PD������!�dYm�C"���v��C�};����R7ߥ���%�
�\���+cSm�n�>��+v	I��%��ik��m�-pwmv�.�Z�}C;��H�	���\����@y��<�_T�h0�I����G�k�$��6�z�b쨴�n(�;ܑ��:�]�O���k;�����GϽB>Ȅ�zj�
cLB_��_T�`z��qө�P��5���؆cd��u��8��] ����2牓���'j�C���9o}e��
ذ�2Ss|ޜڷ�4������4�����e�#K��DS�傦�K�]�K߀�B���&�Lu���5�9uP�O��Ow|�"�ؠ�������F���{z��;g�-]�6���j��j~ד�t	d*NH��g�J���_CyPb��/=dk�w���ɦ�H�)'�_ l2�D�{X��kd��2Yt���}n��~��V�j}��{�0�'�'1N#�!��z$IR�,}w��4�]VQ�� 2u>+Bϛ+���A�kH�&�<��Y���L��2�BL*�2�=�OT�<��9���f�-Bq����g�m&�j���m�}_�^}���e�˩FރJ��EZ�Gi��*��=����n9�tc�=��\���OÃ�Ɔ\B�Al���@�:��p]��WP��n>f�dԊQLX)�#��p ̮S�\�p>��4x�6�;? ��H�A�i��a��􈆆�Û1��g�B�u	M�)�5�������|L�Wd�B<�S"�VܜW�����τ�����O����;>qH��׸xa�{&7�l�v�^�	Z�Ӵ;`p�x�N�	�^�)�;#`g�<4ܗ.�.v���T�-F��m��e�{%*�6K5���i���U�͂Ƕ�]כ�r3���g)�|@:+̔����F]��7���N_o�`�0�r%+>H= ��
p�K☴+���F���� �k�7��QҐN�9YB�s�݀lh�E퀃����R��� �M���~b��6�{���
3���'��1]ӯI�h/Q<�-��_��K�&y��
15bC�GQ�ep�q��������dܭ�Z�h�ԩ�����46��x^:Z����dt�x^�J;�Ζ��s/�-���%�++'�PUO䢬�|}���w��h�\KD���fOG}��0���T�V��P�^v뱒('�ݡ�<:wW��Ff���{�Ab�'�1ѝ��g�`��{�l='�X�G)OE����@��o��o�He�俬�'$,��R������Q��zj���P��6"J\��&w�sdɄ���MI@̐�U��3A T6,k���`�Y��c8Y&s4�"{�&}8qg���ﯛ��9��!�����o��=�!���d i�O$��\��"g~L���. NHIFXo�5�~X@E�����4��'GҢ[����fS�x�˿���q�!�(?�����t����\<�u/_Ɛ7�D�/r�HV {pD�h��K��&[�wH���f���;u�>����]T�����22:;�o���q�
~r9 ��K��m�E��P��e�7.�Tz
���I���E��˜�ڍX�����-��j�:�����(��T��0?��?>��%���h�ܴ-�J�<e�(��6��yҴ��xp��F"�!�}��RoJ:��z��U��#v"�9.�%D�1����F+�D��jA
.���j$���W�����*��0� �ɽU!<�_0���V�b�Ł�F�Zs[>m��m-�����x��4�kf-��Cqc��Lh����D�r������� M9��6�W��NK��s�<�굝g�W�u�j��:6pH8*"�"J���LWcK�oöZ�B����ܰnR�zy���~W�ȪR��t��A8X`����~G�Vm�O��n�,�� SE^���4�4���ԙ�t7c�p%w)��eŚG�u��3�G�&7�A'���I'� ���<�a�f�%WxY�f�����Z����r�*��>#0I��9�p�k��!�9v�����2c]�Bj��'���)[��UN��l�LE����r�1�B=���#r5���[�X�O�3�?�/�*��B���Y��f�9&_�$�b����� Q�E�8l�o���!�H܌s��x�O�g�ʯ(_��l��u�4��M��!1���iP�����t_��P��K/yA�Ovq�8`k8e|vj�Ek��;���x��!8�p�H`��+o�SK����I��A9c��c�[���Ƭ��НZO0�]�Z��{p�g�9�1~��c�'�}�[n�����C������J)(���ғg�uKg�^�t,/��_�n�{���	�&�%�W3�,'-ˮb�a?p4ǟP�)��P~��D�$�dvB�N˒����@�{�1��/~�J1�m�Z�_`�\(�Ha��O"�a��{w �����^s͇�' ���;'0f9�����a��ϥ�q�A�8c>w?���e_�lq+T�]��;IC_�W���,���J�u�XҜ�߅�-
	�}-t��<jxl�[��x�N
k��M���_�w���8���q=����P鴟�&6��	�J
���DL�@�#����快�lZ���y�΀��h�:��,Vi�[�Rv�}�TxCԷ\�aO�MZ�䯩��z��.���g�#r��/�r�i��+f?l�bBvry�8����b�O�5���a����x%^�R� �Ճ�t��(U�)PKl������]����yv6��H��$��_�9u��/�e��^��e�MM��N�����r\�2Q�!+!v���"��;�ʮ:�W'���3���Ee�M��ړ�����'뛇��^+���ݱ������-�r�o�|���(��qU��;V���!LQu���N`��N:5����I!�wH��
�����C5? mM������4����%M�ķ�c֖i��K,&�vgE�y�|�y�N��֡d��>TK��&�[-b5��z&!�%B1�P^(Z����7P�J!Ӫ�IvG������#<���H��6��m�{�WY���o���צ��_!�V ����~���U�s�]ae��>�'�#!GH��ς����?��/[���p��W×*,~'��Zˇ
 ��ѻ�~
\����4ȳsS]�c���V��]:>ɪ9�0�sĺ� '����u3�2�P3>�]��}�A�����48X���|�p�2�)��#kA�[dŏeue�-~?0w�Tx���v��Cc�k�{���~3T/�qs�@v�+ �c���,��G��e��N7�G �Ƹpw�8�1됐E,���Km�3ĵ��
d�{�\J�<_Hi����u�:�vY��'�G\$��S�I�ٲ>�Wp�ޟ&�yNe�]ET�<�m�0�9Ear�Jn�
�@�>��`Zmty?	��S�yw|}�a��˥N�\6���#�;�L���Z�����QF�O/ʢ�t����~�7jG�4���4�GΫ;����k�нX"��e����Bq�6dπ��J +�	r�N��`�8��N�K���v%�<���GV�c����id�� �'�ᔘ:�:ꄶ�m��pҶ��M�n\V%���|*<K��H}�m'��O�광��5{��bm�>��8pfR�(@����
z�Ԕ�K��+�5������M�I2�ŵ->[�wG���k)]�FIX��V�)��ˀ��b�~n�	�I���ώ��_I{w�qW���vB��0�z�f��9o+���GZ�-!�=�IYWc����T�s�'�v���J�O���b6ě���3u����J����{�_�3UP(�J_��0�&_�5I�/��d�ff�g��[���6��}��F{N��v����kC�>����n�q��/4��}x~�_��R0��I���k��ItB��kd����Y|�3����u���X����e�䗫Bk��t��������XJբ9ᶋ�&?mq&p�S&�6w��T�PlަƝh-�(3�d�={8�Ky���>_��Q��YM�O��?���7��*�_��xm�&!���SL%�&3k6��P���(��9u����Hn�ƆEL��QQl�r��.���3�6:r��@Ҋ'p����@B׿24%���[���n��[��Q�t<p�.ă��0�l�֧A)���ڂ��pB�W�p���OswxX��eP]�[��8?�1u�5��}m�+��""��5^^w[װ<)�{��'����g�ŪXR'$��,_2�i��":�y��&)T��m���P�z3=L��j�r�N�ff��k�W�Z;}k��ki:�3�������C�/��C��KB�@u~@�~;��]���A�r)QA�K���>�]��"��Ln ȼ�F���8�����9�E����,]E߿��Q�R��6��_=a"P5���vA�go�Q��\ܖi�?�x~��W�PO8R�B��/A��%%�bS��t�UV�aW�f�B0ۻ��_ �a���4I����N��X��D��B6�*�����I2H�"�J-V�>�WJ'���d���?\c�S̯ :���Dm�%��$	�}���H�>�oQ�gZ�e������>�y�^;5�ƿN�2$��2e��4s�����8+��}��]�K�:M�h�T�1H��m�h�r�-�����д1���8�m�F�H��3���
�ۈ&�wj����3�����E+�hʩLl.s�Xz��	�F����Nۃ�Vy*��V�>\�����aB��|ZH�s;��Ǆ N[M,��a�%�8�2�W3fklN�'?�-.������[_�`y�5Bg���1o;�P��9Ъ4�Ėr��I]���dѡt!rG��[���]?TV�E@�_�F��Z���(ȧ�suD�L�� <`%�	�-�.ȃ�V&�ܞ���0�f�V
e��{���J��/�in��KM�:k���L2�;F�af���ht�,0�P@�z!X���*y��<�䤍h��N�k��PoN�<�"V�E�&��*Z��P�z��N����-��{֌7cؙЋ墐[�d};��і�/��w��ʠ��T�F�X�X�R����.���٤�Ԥ@�ą�5��u�4��6��ۨ[C�U�Cx�h�d��X��������b%�cى���[��#즡P�$ـ�7?� �x\�w�G���߅3���^]���~0#����0o*'Rc��J�$1��{��Y�p���x�T���!���H�x��b;)잰��Π��-�����\?��f'L���IE%"�M8:�R�b�dr0-l5�^�t��'�7NC��cb�ЄJیZ�\��6Ea��mW�!|X"Љ�u�}�:��.]Z��3NS-tQ�� 5����I��V(�k� RuRU
X^˱���ϯ�ɑ��:�j:��L����Rл�o���9V
r3��U�{�D�܉�B%�tf-u��x�[g����#)���u͛"O��U*�p2����~e��Vuh�A������4:"me{N��-6ژ��D������R?���!�n�m���9޸�o�~���~�3�&r+�Ă�N.�r������T�>����K��ZDtk$j�S�(���ߩ�\��l��<c̤w��d����"%ʸ=�����)�����4�Xm�e�ҏ��^��OV^s�`K�ѳ�Ё͐���N ��i`�lC���{��2�.���n�.1N�Ť����z��+`�z���$7��:�"n�ײqU���7t[4�������Q<FQ̒�����oO�ҟ��QŜE�TY8�9���8�,%�<���\��ȱQԀ��@�i��`_A�TtmG�����?t�ax
�9c5��#=��gj��T,ٛ|_a{�姦�B]ީ�Y5���h�m���NpK��G���j��A��]NxtO�!�^�g*�!���8!���G����ˈn�$Ѫ [�jchsX,����,�˃_9��A֪W�F�>�]ZˈD�� *u��}��� P;��p�6L��1��}vٴi����Ga�����Ć�Eވܯn�N����r/ ��f|�c�j��wŀ�r��)�5yΐO���ac�z)�!>.�<�I�E~hMY���ނ�SHQc5&`�Y^凊�!U�#F�q��k�;�g��l���Z���6/i]�M�����j�����Dw�.���Z�_2��#�-�f.�Y� f\I�¿@V�ʫ�r�\H��rߙ��b�:�K����������UP;�ތ��ß���3o=��i<1aݠ���z_����rh|�� �R�wP?�I'x����
�4��c-���m���;~g�PT�d�Ĺa�kF2CS�6�6��eΟ�U�_fR��8��e��((�Ү����ac�P� o��k �\�Q��<���,�Z{�E��(���e)ڱS�H���F�TV+O5��$�xN�	?A�Q�d	4��5W���rj��mPS�"Q �}>�n]�>2Q�����/".*U6{�O�ܩ�@�3�2�p�����հ�R"Ān+�)��ޥkZFt͂W;�G����nBA��h�����\'�����P3��Rns��Z�Z���I��l�?G�\� .�{<����������e,�F7���z�iY�E&F�����j�۴�
�g�R>c���<�.�y�Kk!�f�$���|�l٠��S"�B�i���@�m�̋��{�iW��M�>������<��2���«�Ne��ɉ�al��/��(�-��_��	��D�Qی��.m�L#E�ywٯͨ��]���F/s�=��e�?QׁUf+�E�JX��Z�]�b����NwF��}P3����u9��%4z��+�C��]�D�u-c������	0�2�|��~}Du	�����̬�r,u��˔�wU�D��)����E�0�������5�(�t�c��w���L��J�1� 1G��tk��O��/�[������5q��Z����$Ԅ/��N%�li�S�+?�g����#�k;�E�#���\�T,M��XIj��+/z��u6�rC�f�T6l*�7��6�P΀��`9��G��^j��q=P�����Vߎ�uB$�z�#>��,�T��[����ܔ���J�R�@�(�s�\�8Z��UT�m����,>�Ǹ�Y9��[��#�r��m��wW[��^�A�\�T�g�-E�]��6�2��8,?�����}��0����S�A_m��,��G:�qNZZ��ip�m6x�����j^:�������4����{����̒��W��w���J�9?:NC�ʴ3㎵Aܜ�Fi�h�8O�ok���VGZ��e���<�c�i���w�G�1;Ca�d��|���F�K�h,M6�)����ZwN�����vݾ�y;�N����;S���BV�0M�)��C����P�i�&�<�M��kIt�����_�[�����:4�!af-�����
���Yy
��[W3�ӌ�#��a��L�8��fJ:�t���ߗxEOy��E����{������"���t�lb2��C���"�P��GT.��Nky"����16��|��K�bF�-@�3��]yw�i �$&+ j��>١�x�K#��?T�NT�{��Lh�xe��j�N��<���i���ъ�[�J�ʛj���L ��I�������.�����]�Xڳ1Q,�M.��b�2�'I�W ��
��9�e\Y�E;���u}���hi׵��Gl�U�Q�YU�)�Pf}8|;����}�2	��G�OY�FZ����wq.��6�P�����E�L��A�w���_c��P2�"ދ㹍����A��7�)p�����1;��׾�Pr�����C4��`�a��1������TC�Jq�{(N�vӧ]I�W��0�3b��j�b�i%���n3�A~o�ߥ�O�H�w�x��P��2�ց�|�Ŋ{߽N��qm��$�ri�N���#�+J�F=	�V�������y�U1�s-�-��5{��{6[�qaB�A�M�u]�	k��g�����ճښ�,���gզ�Ӝ�6�SM�$q��|@��&>)�*£���nn�f͵�M9K��K���v�d<�#��&�ח�I=g��*�i��-k��E��b�؉n��oT�wzdIVY�^}�T�]��� ��p�ֶP	�O-�$��|DJ�O`�S��*Bq�;���s�ukN������J�ty`?��VA�gdV�d�gs'�]�d
t��}�%_��YE/�����)�T^%o��)�M��ɽksN���G��=@�t�{�{�ps+�p�����B>��r]��}Ψt7b����U����PMsQ?`偶^��j)��>"u1)�*��:��um�	��01��#��z%��Q|�H�d��ω`vC4j���፿��\{�__F��S��/�)MܿO�ZC��@@����wN!R C��1��IC�k�
O�?00�&v}�G2�����&g�ǈ.m~t�H�k����1�d+UsQ�VI��N��_���I��?�P�K:)���**��9f�.S�
�J.Ц���:!ɒ@�������-��4�:l����Z)"W����h��F��1�A����n��+���6CA,)t�̬h�&����,xW��ڔ��<٦Gڍ͊��#i��h� k~��7��9rl����S�oFb�����G�l�k
�Y��kdf
���x"�,�E�G��#�����(�&AH�qk;YT-��6�^�B�$�/�1�'&�Bs�f5Y�+Գ��-��V{h(��
�?����нb6˜*'��C��F��Aqo��#bYM�x����0n��3ŏKG����@0<�f;md!�v߹2�ِn$������7��#�<�D�tD��%��4MU���+�1DU}
A���O�"�C��q;B�f<��I������`M�����4?S��AL� �3_<,��-��O����M|�GyK�o�^|m%�TB�_��67�E��^N2�<�sD�o�T*��ۛ���������=�K��0N���O�zi	�qM�XM2�
��te1-�`�����:c@��K[�*@ܽ)Z�u����]�X�O+\-Pd��9G)�B��¶����&�LZ��bnU��E����S���+j~��|}o�w�)ie��zrc��W�?]ˤ��/���(W�es��N�9�c58Wj:��Dr�N���V�"��he���Ih)�S`:��lg���fQ�'?�<�z��<;ʈs�������4|wh)���sua��i�^k�����M2���奊�x��R����m.A�z�������y	��n��S&�DA���R��	��۝L���p5����5���&#&���e�fK0� �Ȥ�,�̢��� �[�?�w�<ȅ D��HC:B���,h��uN��O~��1�5���,�H����\��khS�� ���D�
�?I��gؕT���	.�]�ъ�P�����?79��������9C�z��޼�S���P¥}�Xw�2 �cB{s��?�&�,�)��H���P�0F�-�ި"�K 'f�@���ݽ��o;�.��5��L���g1�z�3B�������r��>_�����(�<L�|��46JM�)2l�K���:�W{����p�V���ͳ8E��2^�7���t~M"d��ET7�+-�Q�BK�aT�*��� �Ǯ�~��B�t{����1����1���� �C�~� �ToaD�m-�ab�o���e<¨�W#V7sxa��:��)�X��h"(iFu&O[�%9G����h���T]���b�WX�lC+��+^=�� {���W"��P4��"ErvQH�[�I�Ŗ�Nh�1$�6L�!�[:e��4M?bM*�.�;-��~�_r�!>݋Ҹ�!ޱ���@��m�zJ&K.����p�ˊ	��%b��)�vu0�@�RK�v�s���C�VA0p��T&ȑFqֺ�q)2�l��t��]�|Bt*:q�$��0���u�;#��-�8�$��2�S6;�D6)ǂ���WG%�*�d�L�G�Ρw�&����6u=`<[R��Fߟ.���L��cľ�U?a��sG9 �k`����r����u�2"���AY=r�8:X�ͣ���Zi_Mj��N�bFP
�p)���+֜�-�?)RP�82E	e2�X/��	 ��i��m�k����A�J+}/AW���Cc�]�ۙ�&)�YfP^k����"��\�Y��T.C��O<=�ߴ��}(�Xa��zX�@6M��hF|��VZ�����!�پ(���%�mw�_��Q-���w{Cg�����O��_;��r�e�O���5�&9�c�g�Qy�j*/����&��'�^#7�r��UzBw�Y�dV�������DF����kB��<+��A*�Y�ǥ�9���	��E��O��W�����ڗ(09F*O�Wl��Z���������S<enl[	&�F�a����H��|��mè,}���1������[è��Q���Ak"����
��(w６r�擝��Y��� y��8Sv~^Ah^��:Վ��]�v�]�to��Z`���zE�7<�J��z�����t���fa���t����JP�D�$�
F�v�
T�4�(��BC=�M��`ؖw�UJ���&�l<(G���IsG��xtaq':�����G�e`�
@�M)���{�"�Uo�����'&z���J� `w!�2A�����q.z��n�W8n�@����d���O�G�����w���H�&Έj����R��Js����	WyR�=�WӱS�3������,i�x(��@��r�5q���N;�1�e�X"�-�jH���+/��� f�ږv�&RG���$i�!m��9����Z7��R?�z�z�uͻn��H[1W��6@�m�ꝵQ5�(���C��~D毣�"�����N,��+ZD����;�
/�KM�\�D�c'#=3.�I��5w�W٢Vf�~;7��o�S: L�G�=�rr�����V��H��T���?u�S�l�J.D.�R��б��
x�#��usD���ߓ>���sl7?y�W"K�4G����8��S^��p�ɻf���6�U`���нN-��c��ab�S`L��7>:��<:�4]Jq_�R$��,%��RO�RR�B������x�1:]��W��at$9*h��-_�	o��YNJ<��W��D綠.��꽙�
�4-\�v�K_m��ps#���o�ԉ�~�6m�Ș�Q��?�B)���R����H�%�G�O~��;�b8ӌ�\ja�0�0Q�Ъ�@�Ϳ���Ew���Q(R���è~Vz�x��T����2�;�x_⪒]%��҅3Ws����~W���;G�~4ΉN���NX���W��N����jkeaw��������cmnV,�z+a�$|��mjT�I6�ܱ	��Sx� ��
:�D<�<�O[�E�~�6a�F}�����ek\H����>���;Z�	�����;��1��������4���v, �"���l��-Eq�,�!�I�X�u���n�=�S{n���#9i�� 7��v�p��q���qL�u7��U��P�㰧&�����&�Mw#ŜgS�� ��V�AoL8�FX�I@>Q/��Xا��_6SZ�-匧�w��}�!0ҽ�0]h4�J��*���#��[��T�%��Մ��X+��"���ƀPXZ�����p2��Ă�-��>�ho/�cK�ʻ�q��x?	�f��
�]�
�W���A<_g�xQ	���U}h\B�{4G'���O=]i�$�����%7t��T6(
���f��c��A��7u[:��>�c���>pw�\[��'}T��ǃ���Yx��S����K�S��h^�C� �7�()������,`��ϱ5�\��q���`
�˷�;ꗉ�c:w�h���n�B���Hd��`�ZD�����i^�Rw?�=�{9���d�/��ػ˯?��R�z��>-�%�ImҚ�a���ye�y�Mx��^�X�j��N��H����2[�GU��pן�]ۨ�}�?C�.hr��BI*|�\��m��ѥ+�\��Q��dS�Sm ����[��L����:�\��9�]��x�Z�]g_��ܥ����6L���_b�h�^��i��A=�"�w�<�L8ѝ�Qe۬6<��L��e��ni�	�,@R��5��^Z�e��[CP�9,���H���+>���DZj��4�3����3�ӮQ��b?��rˋ�G�)�I����۹����!�t�ڨ>�L�����������o�+�ȮD.y�����-�ZTA���t������<TC:�B�t��:���pE�M���H�FnV�,���6C�������#�'�T6�/ޒ�Nƍ��-7�I�uRW�3���h�ۚB# ��6(��)��3U
��Q7Y�b�0��h�"���Ʊ��7�~����b��0�ܟ�����QEy@�W��J��))�=�TK!��]<㙮��1MSW��r:rj���>��"w�޾W^Dȭ��^u ��Bo׉�=M"n�� ��'ήPQ����1F½�=C+�m�ݦ��&2/�o�@�t��m�t������S�jn�*�����%�����0����d����-LvOur�W�;���jE>w�����9k4�1T*,C�ZH��1ġ������d24�NU���c���@?�Ûr��ur�B���\���NH8�z)%RM[TR�����-g>�kC�B��XIag{]��PW�C,e��uE��͡��]txz�<L���*�)��F�Yu���C;B:��8�m�P�S}d�����(�950ҏ�9*��V�m��8�u?|p�kL�A�K��ߪ@�ܰ��W�1Rj����q����=�%�ü N\@����I��ߕ/�V:r�࿯@u(�j1��D���Z����	G`&���"�F�Q��;���գ1�I~�>��8Y�/����f��j�X�L��@V�%+߽Q*� a��z�&nǯ�X�'�f,���1�(ܸ�#]����,א��D#K�s�](��іA����q��!a�)ѥ&����?��#��\Vr�9�a�k�w��q���	�[����Ѫ���W�8\�2rVd�O�	{
�=o$(x# �e.u�,�ϛ��u���A>_�`��Z\@��cԄ�$���A���`�s���i��H\}.���F57,iE+3P�����Ԩ.u�{-6MQU��0t����J�Q��S8��:'�*�ܤB��K��+��⡚Zi�y�JȘ}�k,e�u:3?S?o]t�7+r�Fɱ"�4�3�&[�gu�p��e�@6m�+ڱ��������.y�5*<#�T��ٰy�|Q�:F���i����%o=	w\���f8���<rj�pE�w��)�yF���Z�/ lì��%��u9t�@ˢk	��� p^�5,5�
�,J�]�9xiaM��f6�]P��2�����#��`���[�K-r�:l�xUd�X�����g2g��z蝘vM�l>�|����5sO��@M�s�<Ḣ�}�
��������K��e�/���+������"Z����K.J ;�N��o?r���: R�kT��� ֖)�|x!M��q��\�#�ǽ�V�]꿬�)�y8�ϱ�U�`V�3�hˤ3�׋}Akcn��*�$o���e���\}��9���'���dv��kV��|��/QNK�=|����U�S���Ɇ��2A(����V#���#(OH�O0��V�e����e�m�W�f�}=��UQK��5%��	���B��mx��Tl=��HҮo��!�i�*K�	h?���/��ɥ4�<�3�p��,Ζ�Ʉ��r��tO�l�����'��@q�]�[�������y��UYh!
;}�k�nkw��44��dۨ���5�	�J��h"�����l�e�oF;]t�<� GtS?(�Z��ERǷh�[�ɕ��<~��Ji�%�TW�¿	6�g��������d	_A�)*ƴ
�h���pY���s��V�u��	e���W�����[�0z/�V�b��ܢE�Q��G���5x�)�������}��	o�u�����c�h[ rܡ��Z,����V��^����W��q9ٵI�,z��O%�p-���6Z�f���-x��Yn��~�@��C:��_~�YvjZ���X���V�0��L.|�#�Xrʆ� �%]+���!��R����ԑ`���ީ�ݑ��9�N����m���e�)�m�3a�s)�$���ng>�z����%(������ג"����d��]���E8����@?�Ⴎ�xC��+���Y�Fz]��=0h�헭Q��Z�2d���Gl��48L�[~8<�%֑�����ߋt��ƐJ��8��_3�����&��}�@0j>�!��Eu���!_D���*��i�5��Xa�z�d��n��e��'�P�Z48��E���;,�>�-ʹ�ɫG|H�Ȯ<� 9�s�ݧ�+��лW�
�c���J�O2��$�D!j�?@h�^{� �8-��0Ʊ|�6�a�S?�����mc����x6�)�&N"z㰆�1v�����)��b\�0�h��m�<S���\!
��h��1�UaS�zwj��z�r���X}%܈]�vu�|�ã�jb�����6rY��W�u$�D���\d�_�s	�������HJ�w�`�7�]I�,ģ,ƻm%hr�y��N� ��G��D*�#��/$�U$
�A�81�g�n;Q�mQ����[�)ܤ02%>� ���P�gz���wQdC���%Tn��TosF=@�I�G8)+ѽp'��� ND��<|��C�_��N\�U<`Z9�d��@��vQ����f3�҅���*����o �\��I�xOw;R�֚dWn��L��*;Vc�!hG�y6�c�E�t��N�vF��K�0�r����ʊ�9&���ee�������w��j���k�����"����9��W1�E`�ͭ?'��d�'[P�����]U#�ĒL����?�2X��d�=X{ݭ�`$ν����B%)����୐g��J���Jڄy�ȅ��Y\���-����c|>7�8�d�Q]�������<��՞�(��A���.����ɵOEJ�p-55�{7��m�8$J�G3�`L�sL;����W�[��x���@<�+�Gϫc�Q`E-��m�wWb�K�1-����B���� ��B��F�ȞiC1P���dɟ�7�AǑ��G~#;�U����_C���ￓf�����]������L�D\�*�(�Z��al�!r�i��L^A7�0�1mwH�k�N���ѡ�Ɉc�����{=�~������)e^]$�D{7���_��x�/P�ٲz��F���g�֡fe��-nGz�e '��3�0�Y�b�����~�7h.�����������cF0H�߆�!�?���'ڵ�)0��
���ݤI̲X�T�9I����R!����vh;��(��y[�d��WN��������l����Xk�@�ݫ�e�����(��]�	J��&�y�Y�m,)-C!�!r���:^�b6���h7�
z��2"�+T�
u�svR����Ǉ�+c�	{YA�g���AH ��gi&�)Ec�<��1ڝt����Ѭ�SX}2q�ɭ���vMX�]]�RJw`�������H�sxnG��W��6�X}w�4]�Z�&D"��#N��=�<Y7#
aC�)�89NSPRj��
��	�+DX���~���aU�TV�M�.�e
��v��v>�%�������8�%�B9&�8[; ��%UZyO�M�X~�־V	�:�h����P���c{]��N�C�OO�[�E��lX9l�P�3��`�wέ���z �*�Q4�{�����Nd&���
z�������ߍ&cD��f��J�vt,���Kf��dہ2���UE�CI���+�	Bu�7���D2�c��k��`n�牻'�~��c)�J���J�G�I��ܱ���礔�QP��	[��ii��;�j��z:+S��Odn������-��ױ�����҆c��~LN=^`Հ�g+hJ���Y[�*�XS�0u�g!X��ӿ�v�P&;��qj�zH�8�
��)�^/�5�tE�h*���2�ƁxN�M\M�Z$�U�(��d�:�01�0VOμrk2�g��֙��7��xg���,p��X!��7���S�C�O=f���E�R����N���{l��毣�&�I&2���'����2k�d��q�V+T:��z)��^�LWq��Q�~����is�s&%�p����Bƥ9������`�@��v���p���K��V��	Sf�ԥ��X��m/�*�5s�Ћ��aoW�S43�J���0`��>������s�����O�酕����G�\#�_��F����v�\Κ�`���I�`V+;jM��%L�4��gr���f�Ć7rY�NO#�H_�9���S�9������U��б�ɉ`ZG}�]}��Ig҂���T8��z���#�yw� �?�W{�.�~�+@�ٟ�����}��}�R57ZXPn�>��,������:��uy�i,qm��vyr���h(����q��h�=v$��e��|�^,c�~U�����fқ
$�`l�q��N��x����Ј������H��ء�;���jF�\�UtA�!dJE��\Br���>��i���N���>z�ޒ�ӣf�RR�Ilg�O�.q�@HU3jN��c�lϕ�%g\��e?9�~r:>��m�9z����q��P�(��QnȠ� D���s^ےaK	I���=>��.��v�����N��BD����t�9�����s�(�'
@
R·Q$�k�Y�M�n)�dV�۱����i�!I�]ډ�_����Z���z�	���?{����Oa�>�'(u`�V ������v�߀��;���1��냠�|���2s�~��f?l�=�����;��%�v��O�Y�Ù�����B.��>��$����G��P������=j�[	����$`�r�X�c�s�	}"8
��J�jQ��X��hn���Ȅp[�,�8�s�9(��$@e�Z�48l�,]���!�9�~\�,"=]���O���ꪛUi"d��2B�`�>1�E]y��G���4��X
v��6�`;�G����*L�B���ǔ; 1��my�-�gl��k�׵m�^Լ��Vìf��1Yػ�9��J����h�-�6�����h�<dgC�G.xbFJ�g�� ��������}�&N�o�ӕo�k�z�6�~��W��W��c�\���X5D\�	�;��6Rb�+	�8xϾ�8E�Z^�������.; c�:Q}=)P�@�]C!�a����O������P�s{��F��ӑ��Ύ(�v}�;x*����e��"���$7hI֟��9B,���E�y����)�|�<>�����ĻY�D {dO�����g�Il��lqF����$�4��|*�.M�� ��%lō�|ȍ���)oODD�����x-���7+�j��U�T�V
����xg�v��ʽi}��� ������ө�S��c{���ٍ�f�M`�~A���#������V+	�Dw.�O�id�)`Ҝ�bZpti@$j���4���M��h x�;�#oX��z�MO�"��^;�Fn��^�������L�L�-�enz\�Oe��`b�٠ދb=��̸_T��C�°�s��������E�����»���QY�j�9n�A��f�k�,�"��.��\��a�z�GJ�R}@�Z���C� ؐ�T�9�dѮ�@ V�Z�ȕ�-o�s�9����6t)6����(�`�lGp�${���_1���F����8�{R���?B�u�RAZp��b�UJgm")�:��K�WǑ��)���+���y����?���2�&�D}4��ė��^O��9L�!��5�W���|A@�^�a<�!��>}�~��?���yי��r���n2d������"�v���p�q�]�Q��G �����Z�Z�x��a�o�s��������#~�w��H�,����f &����U �  �;�إú�+eG;E�'�?±�|(3��	y�3�H��tVz��e�$},���.djg?`I`!�P��M�Qha�I�+X;:�]}\�J��X�Mh�ţ�,�`a��l� ��ǑaN,tyk��+����{��P!����GM�0q_E���1	��A�1bl��X���C����2-�0������*�2�8}-s�[�u,Tb~�!3eE�
ݎ̓�#��h�������[rbL�c0R|U���P�svEE�k�N�*�.���	La�('�jf���?6�0���7h��8Z�`-67ea๳���0]��x�I׍��Y�*��U����nw��������ԅ�Κ�Ѳ��|8�kn�Gp�\���̋�`(�Aޏ-�,y���v��m�h=
x�x��@5���	�X@��VTQ�a��x)���1<���������/���w�_���V&pK&,j��΁9��1(�w��mf�ԥ�����;�}D���͍�b#���:&L��Uz.J0-BpV�#�5�a�B�'I�v[XK(qږ���%"�M�#�]���N[4���{Աwh��)�0���?g�k+�����/����.�-i�4u:X����rl����]ѓ�6(M�U�/7|���3d��%� ���&6�yA�5���y�ZBT���2���}�����[�B�*�괤��Y�6�ߜ��<�������a�o��� �.QӔ��W�b�����x��D#ܖ���nQ�+��3��!�V?����x�#qS�I�L��Ѧ�8r���^ͥ���u1(�������i�����ҝ�u���^��7���hx�b^�����G�Բr�TK>"���:C�ĩiv�#�6�SS���ܴF��K����Ċ�ڭ �q1[���u7����M�C�g����\�'i�W-��� �ናщ�N��S�B0 ݁1�s�:Dv��!������cm���]�x��u��1Q��>�Q�2�p�y�|\T�`ӗm݋/s�.:v�w�N��o]��{/�(�.T�l��˾��믎����� 6SS�����<����y�_�t�i���BÇ<J*����M�!����û#���8x��puӆ�V�^�� �y�����s�^p��I?�k�xAi �� 4L�U�7�ܫ5���-��H���d`k��7�$v^����1��/�A��`�2��4C^�Wu��@)!�,e��������e��x��zv�.��ϏBQ����U��Ϭ��>[�>�:�i����D�=W3�ٷ"K>�J[�sJ�)B�}{:�M��[=�t>���zm��4�S�&�%>CO4�ߋGa_e�8w؞i;��ʝ�����I7���x�js��/�2`D�64�������+�6���r�O��9�|?'��q���ǋ�q�Έ����l���ܛj܁4��HX�#Ϝ�U�GO�-�1+�~��,�g��LjZRD����ȅ�P��`_��P��"�ɮ>�o�e����}1da�P��]m/�a"�����E�7iU
Z�T��g�&(0��� 2�b7%r�K:�Ȳ�'�!.��yX��Q�6��_I�$)�Z�w
�;�2�Д�1l��c5:�4ʇX�R��7���7]�C�x���%���!o=�5��~�2�B��w��_h�wU��~T�|&�Ӻ4�z�^�rnݐ!̲Q���-���� ��MPH�ï(
�J�,��75�'��6�?	���Y�s��\ׄΙ*E��*�[���A>G�.��m2҆~��q�"p�2q:u��!�U9��ғߡ�����g��9�uk�.E��59�}��"�C�����\gw`��\@��������ʥ��F!��NF�cՎ��4���K�����n�T#ւ��Iyr��v�C*�H$K�0�QN��p��ꗨe�l�)�Y�KǬ�S:�����\������10 j���%�|�����C�B'&��󞷩dRh��di8&�4�E�C>��G咖����h��H���y2&v�JE�sJQ��p��Vҙ�V&d��B�*<���]>x�}�i�:�=�m�&C���V,NO�y�a�A����6�p��-u:d����7�e���-�;���R~ ���+������s��k3��ˌ��>6���p
ο`|��Y��a�*�+����D������}�O�t
��B]��E#plZO��퇢�z_Pc�=MKw�.Ͽ��.����٪�cݜqvW�5���|�֙cX_�1w��E���!�V낇=�c�3�������х�!���\��G�W�@��8Y3�!O5�L��\rC-��n��ި�B���ƊG��~%@Y�!�[焱ֵ�� p>��:�h�VwiR�"R�C�޷��>��=����Q��ۿ%�8�}���z'k����Fss��29�l�|[`ݐ�W�]�f��AKK��B������6�pƫh;9�G}��&.�ʸf�1e�Nv]=&�������ӆ8�-�F�<�񚘤6%��7��CD��1�朞��i������B��)���Zۗ8���DG{|��\�B,'���X"T_�u�뜍�)M�6��U��PM�nADD��.����RyQ�N���d*e1�!�'06�) �°������7���� K.� ��j����e��	��- 
x���`�	L%�Y�`�|���r�FGW����,��S��F�N�if2v����in~`�]ap	�ݗ\^����v��:�-���?}%��W�pe�GQ(�n��lcG(F>x��R��h����R�K4X�&������W'��G�<z��w��A|LyN���u ky�g8]IRd�Iϰ��/�q�!��ƟH��-\�1��
Z�6[hN�E}Xۼ�XIO�>ɪx'���b�nρ)��=3)@U��b�F�ӛ�D��\���v�Hz3���i+��x&}	3:!�L�YT��Q��s�i��/��m�;_1�Q�V�rB3�W�O���۹<nA��,mB���&�������̈́6�6=5Bq���%đdê�V��#�ٍkf��s��� +Q�8���nF��WU�����h�F�@�i�=.�{�(�&E+$4�Nh �U��5O	5��YR��\�r�����lc���=}W�S�������
��y���_&ۂ��m���b���4��um��;�?�Z2O���Mz����;�$�+��C�T�͜�MT��d�8���g�o�4���o��-�M�i��5R�m�r5S Ǧ��x�����չ��G�����,vd�q"-vT�:-qW��*B���w����46�R�L{�Q]=o��v�
~�������N����A��^	��KT�(�����Wm!"�ΰ������	����ׇ!ѹa�.�i� ���I�;����\�ĳ����B]m��mt
4X�Gfca0���.ul��-�p�ŵk�����G��8��>��-i("P����u���<��~�h%���b��H���';#O�7 8&��oG敐eŏHp�6g�I�t"Ū�?҈��_�["���a��rlz�����=H"�wr'+�.�a�E��Hyg��J�_����(�sw
��X��K�Ӿ���`�������a�[#k������趾��x��yw�����/�ņ��ۧ �ӛƣ�����Z�<��MgBA���P9|k��	T���w��R�K��'�p���v^ �x��R	��&��@Js��Da��0�
 B�lW��(b�%�i���Z���&�-��K9�H YMu��~�Q�J�o�Q�����YZ�Vs�Y��$5��i���I�����w�w�"E?8��y"=N�̓]+��i�x7 ��g�z��#��v�B4����sr�����Q%��P�k�%���"�ǣ@��H{�B�	��Ø�-�����K�<�wlw{�)*�Zr���T�sĀ ���&1K�l)��[�q߭�z��@*�*o?�A\C�o�{=���`��zb�����R��٪{2L���q���3��(bX��`�b�ݜ��z�.R��/��	�)��⢂\��}�w��`��J��\q��G˒P�ʻ}��&\�#m�Ѷ6��X5�H�{�ܗ2�Z�n�"��6L0�⇳�Z9�Uv�C�e*����P78y�71�w氌1�xk�T�Gd�%c��s`��^/A%�N��y��`��=�ڽB��O�DĘ�4\߿�����%ۆ��;1�� �t�nd�?ⵂ㞱t�4�%N�aฉ��� �Q��c�#)����q�$�f"�g��6P�J:J��n��cW ��IE.}Y[�E�u���5d$�	b �k	/I��	A���;tw�/�P��qb
��s�6��E�k��4���b
���FY��r0�%��<	7H.�jFY���"�5۔6���ǎ7ɿ$���<�B�s��.Q@CL�.��Xc �����D7x���h�g�`�<X(�=Q�����N�B�f����pB�Z8|S/b��W"���v�u�����c���&|� m�v����S�pGq���.h&E`h���ɹ~F�߮U�fMȨ���%��D=\��x	�7���l�C�Ix%X��X�	}P�u���P�Q�N�U�J�3��8F��+�=,l�i�B}  �&��'��Qq�ˍ��=U�<���}�(�mg�Bm���XAd�c����ߘ���ג]�>Ҡ���e2�{I噋y;�`���z&��hH���h26\�DVO���Q�����u=&�1߬h�����z�)f�e1W嚃�n�v��d��4�ۇiY�����ͪD�8ܲr��DT��[�s�`"�/=pQ���Mr���גfx4��t�l�Ov��}F^���m�tB�'l�5%��"�����O����P&�~��b�����3Gx��;�G�^�c�}��gT�>u���;�[������9�4���Ǖ�4���ϴ��H7���i���@E�6��x��ǭ�'f�P� �b�D���bS��a�K\U��=x"�:�|�8'����3	fƖ]���Rn�s����R�u�F�a�*���2T:֬3�]j�LN�T�т��`�c�հ����ʷ�,��/=�T���b���[�#����ziW!����s*E^�`�*���j��z#Ⓛk��!b������mRdR>�������5^�5���{��_?�n�o��V�p�ێ9�����A��h���٣T)�V/ѫn��%eL�0y?��;��W}es�.E��익¶r�xg��7�e���ɛ<ۢ�=�2: '����+3�W�]�4c��s�Q�n�O�Nwyȉ����ޟ?l�+�l3��8Ӳum��:p[��,j1_��U�v��T5�޷�?�^ÀC�@�����>j%p<3IsɌ��b8����[\~�#y��&CT?�K[�&��K���)m�iu��q��i Q��Y)@є��y��[�F���T�#x�i�|��ocu���MW��?ntFx%+-v�;7C�!��ɾ���I;%م�0��0����l�ѽ����v�trx�LW��5"m��8��:�;�جS]̃�!`��������L�,wMf7��E�f�Q,-!��"�������0�(q���ȎU�Y��� ���b?g���`� #ZP����Z�Mė1�������0+�'�e7h:��l6D&�-t����-qxr�'��J�$h����Ü��`�ڂ��'fG-�U&��	�̎�C�1.��-)>s9�Q�b^���uSpj&I��"�F��L��k.A�,�	��O�x�������)�Yc���<q��e�֚TV�<OԚA,��-*� y���/2�H<�:z�ObϙS�5ZV0𷅚��K #�fS)	��3!6Y���&����h�-�𳬈�wȮM���T]���KDt�� )Li����Z+�W709d(��R/B���>��c��.�������.#ް�Bg\5r����7�*e���`��a:�_��K�O�`/�OT�6��(�dwH�4bĎJ�0\<��C��2�Y�b�B̘���L���̏θ�F��N+��ڿB3J^�|�(q�t6����|?�H����+�g؇�m���U�k��A7zbNY:���C5����Yh������.���v���A׻6�����n���x�Н`��8;dֹ�tSR��G�ꨕ�e����&�2E&x�o��SCm����(N���8s�wG>K����u��>7of�s��]�Tk�2�T�W����v� ���ɭ�kg�w�yh�EkVs���F��q��ּ��h�N�8/=�����@g| A���9I�;����q�tާ����*}��F��r�{X8_�9;*w�b}B�$�U0�H�Rs�,�0Thũ��G�r΂f㉸KI1�e3Hqlo۾�܉�qP|z^Y�m��K���s���e<�ʢC��v��j��nj7�s��F�"��[OxĲ�: ��D�����Y�wA8�`Ҿ@{'}�p��#�� h�;W�ߟ�~l ��5d�b��#��fh
h;Ԩ$��l}|-�bn!�ö�0��"_����3�oRa��=(�U�?�Y���xRR��aݬ;�b��l�6��Z��NO�}B�`��@LK��׀S���i�X���}��=䂏RyKT�����Q��Z�fP�Ϛ>x&Y�R��m���=�B����V�S<��K5GL+Fk`Z��t�Y���s��+z: ���戙������M��v;=�"�]YM�'�����y#ꃯV0�R�<����!1&}D P�_b%w��T��*���	�`k����>x�]�x&��G��q��C�ZeDeY�0f�\ʼ��Y����7Ni���4~�����9���Ȱ��I�n'őa��wy,��#��b��3���~�NH�0�ٚf]�������N|Eħ�+W�;g�U�(%V��/{pȖ��ܚ%�W.ȳon
$��������m�!�,���U5:�w�8�7gu��nF+ɊA3���L���ZZ�xo �ψ1>�F��⬮>h$r?c�����z��I��x��uwj�}Lo]C��kS=�BT�衦z�&��1}7���:�Unb�}����T��l͎d��-�uT3d�j���Ϳ� NU+�̃�L��7��Ah+�\��[7O��J��c3��N(N[�����-=�}
��D0��%�.Rӓ�+U|`6�c� ЉO���o�]+���%���nhH�f���[�Ot�;3�9�R� �Ys�UB�x6A���B��S	�Y=B1�8�<�P:f� ���"���&�9%��R
 (�:
����Vuƍ�`����0#-�!��ߘ4.��D�[ ��ex��`��o��9�qpm�>o׼J�~�Źxϱ�.�4P�ԻѴ%��[����5���[�֖�
�&·@��9��c�g~�O�<*䇧:Wg1$`�),�[�`��R�;����~����w��AJ���GҎo�},9+ �����}��H"{Gw���4Z��镘f#��&����=i-��%�,@u8\�j�,�"��*��{�|=Y�';�"u��1h�܊�'Q��X���F��l�f!&њuZ/���'s���x�hshڏ~��i��[�8t->��BQS�>T��-3�Õ2���Ck��=�llIGdxǻ]Ӎ:�% q�M�E���'�
v�� �5�R�w�J�|.0�1�o�1[TW��C��/��5����o�z�����ց'R�g�j�����)E/�:��Ԝj$��w:\[�&�feBGC�+S嗚�J%}ӱ�ɓW�AS���u�sȥ&�giMj� n)��X`qr�
!hX��*۬޿]dk��PŰ����و��>4(V�!�R��{�V�E.����� �]:
�!Oh��
�<y�u��9�Qs�lqq!���͵��)�!6��������B���ztZ%��d���c����?��@���3ѵe�u���������h�N�m��y#�y��q����3�W$m������ۿ��%#��T�]gL��O�$�G�TB�.8����jHJ��m��ї���4�_���_l�+m~F`��{0,Y�r�Y�g���7���Tz(�r1�cF<���HXz�� ���R����Px�{Å-Z�o̟�J bGFFĹ�YTE����EI�!�3��C��g4�D�Y�#�����v�eY�d!6`�)�6Xޱ�7Z�ѧ#O���TǙ��:o�=;s�}6�	�WL?_{���L5]x2S��6�yR7�gs��c���Z��%�$h{�t��.���� Q�Nfj����ǀ�;�oSO�o�^��|� q(q� �ᦧ����%B��rH��ԯ�u�{?����"K��Q��\1/������2K,:�%�>����
l������!�Ф�g�h��Y��sQ�u�J_5pO�ħ�0����ʂ�� ����s�0g�'޺a����Y�/���tFr��C��C���c"��L��p<��8=	B����Pi��k����M5n0��$�$�r�u�Y���;2�dy�>x����_�l��Ώ�.zf�16�T���,�2]�����W>^6��$6[�B��8��^��.?<���T��O�>�ő�~���?~�-�l�%�Tb)�e�(o���0$V�0��IB�Bqȕ!�<ȫe���/���e�l ������jl9'���z�݊��Z��F���x���� �q֙�B���mJ�eq�p����o�sZ�] qӋtR�T������h� ��0��0K�ci=ٻ�����.�ͯ�d�U�0�% ݍA�²Xг��d��J�Jm�����_�W�O��A<��8d�����E�v�6�����$�o����e_��Iޠ�ò��B�MA"�eBHw*+|�=D]nGQR/��x�!-��}���4���n�LB������	dܽ�SJ�_v�0�k꺺�Y)�G�s��Z��9�3�酈�٫y��7��5���2�ì��
�R����(s5�S�^�S��M��G�ӵ1�8�)$~�ܪ#E~0���?�W<���x�]��ꬭΔa�t���B��������W�M��kLѨ^03��d��q=Z>��w2��7ig���J�b��J!����փ�Ưg����LE���N���gt��~�Ta��:�T#�ҫ��.*����׊MiEǌ�0��m�Ѭ�4i]W�V[��X-�~a������[��4q�@�u�T�v,�����%�l�m�*Uy���X��d��i����n����}����3��y����ڷ;sP3�4�~{�]�u/#V�6��d滛�!o�"5p����#ݪ�\�t)sdv��1�(���o4�i�"��~S�N	-�b��0mG$@VDx����mw��ypSb��DIe�/�5YHz� U@'�R���?_�b0�ᛴZ�V�ŀ�t���{pB_��o�jB��W]�b�l��6�n�Ed�U�Җ�&��t��"~���q�-n q�>O�}=��!qW2/$λ+�cE�[f*������w`��v`��W�,��v�fSՠ�h��PѲdot�<.-�@�C���*T]w�JOQ0yɍ�J#��5��$�G�����A��E�?Um-��h ����Ù: ����u��	���#����&X�l[O�ڀ���_rr�	,?&�;�-s#]����-�V/]���W�&̟�Kȩ��|��A��pFF X�o52ޔ�O��-��l�����A�M�J�,� ���.5�r2�i���frV`ۣ�t
�V���<�����	G���ny�)cH�bľwV�Fl>5�Mϐ-��k����<��CT���%�a��8��m��<'y��f��q44�v-�%�^�F֢jv�,�j��L�EO�O" )-Gn��|�����V�I��+�� u�"�@s�暳���&&�{f�5�(�a�k��
W{���M�M&�+B�S�l�v�"C8����N;�x�'G}8�MM�E�|�,�F�+H��P����9����O���:T�l����>C�]�4kF�c$����H�Z9<@��|�2y<�K�(�R5��p��"������L�%:> u��4�4��C5��ѽN-Jn {�Oz����MNʏ�"�e��l�ӻ`�Es�2�Ao6�?Z�A5����A�#�(�e���#��p���9�-�z�p�
�Ki�UD"��ܭ/�v�'u����z�	�ej\��ԏ.Ъ���ƙ�?^;Z���{J��8�P�~����z�kTt,Z������m�~༶*�����(`�3���:�����~�!�Ai�T�!������O�5 匄Ý���uI���g����$2��A�P >pģ����fF�VA��Q����Cۊ�^>�l�X1��Ì�_wrw�@>)���5�����?Cx��*ɳ����G�Yl���ZG`Ԧ|_��Җ�n̵�[e�<Ôb��DN�8�5f�v�9"��q��7CI�%�F��@ͮN�3�P�G3�+�x����P����p���B��f]0s�5��')�
N�O]���w����q��{�x�j�1+ ͂N�_�|S��8_E{��O����8���%�wx�+�P4���}Dn˽(��J�t$��ˮݳ���Afݨ���O;1��n�jC'�T�u�~���3%[5�!��s�Z���B�����~ߍ���Ag��#g�>e>H-J���F�X^�w��^#n�>z�d�O�H�cra]2b
\b�R-VP�K!�>
�Q�RD@�X���c�1XV���_춨K�S�Rf��g�ȧK���\UCq}� �()���g�! �|d�rD
��^���I#��o���G ,\��y�gn���m�����%'p���w��R�X �_�	�P��f�&�=��U�$��)��	�#D/ԇZʔWgXj^j#�Ҧ���۱�vQ�!1�3:��n2f9��ihD4ln��F���x�6K�G�c:;@`��Z9M�QZ������yC>�T�{)tx�3�)�O�F\���(񅱖�w0��T�jf���jEDf�S"������Ķ�(�fs}0��Z��U'�����m�Κ����z��G���qݒ|&W�x�~�Z�V��H�D�5`"���<�t�r�ݵ�86h��i�$�:��T˴ܴi�+�eBe���e�8�i�SUG�W��`gD��j������w>���[�6d����8E�XT�kj�P�n6��t����/��>H@D.v{-Z\�N���r�(�s﷨�W&�b��$�oY���9������d]�����!��#Y��px|_1&=
̇\�<u�*xy62��2�yD�A�H<��S�_�}�vw�>Fջde��9onE4��'I�,eݺ=<�:�,�OЧj4G��_a�;�7+��Y�p5?	$�z}!�ѴkU%����#�q��#R���.Y.��Po~��5T�� ��'��W��[��:�s�f�2�<G����R��rf�2^w/9Bm��"E�A���ї����8ϰy�z����K�L�1g���v��[�Ȧ�	�,U�����YwXEur톇�(�F _f�/��p�!6xj���)K����=�޷e=��03{���f���
��V0.|�� ���J��XwN僎63����Y�2O'�WD��qy?�����D^���h�{�!XY#"�q��L����c���Ĺ�b<�nq�Ԗhd�����-���e�d5�sk&� �8����j5��-�Q�>E��V�.Z ����� �0���#ڭB@ً����wﾰ�FP���jĝ+�� 8�
��N*B�>5:���u��-�+����r�K0����&e �ʹc���
��%Z����^]Ԕ��y;���Xǝ"����ʛ�?����U8��������ºA):���0���j�tR���AfM3�DI/���N�]y��>�t����\���ʽ���+]�
ӡV�^��T�j6t�>Z ��Mco&n��u��uTbbkS���6VU�Q~�]i���p�/������W��_�7[���}�ϓ��b����2�W�>���r��/ʜ.W�Z�b yJ^M��Y4�)5H��<������2�oJ�����rО���n���u�~@Ym!�X�f%���8;f|���/���Eh&\�e�掰L����n��E�=U��'eA6A�+>ڀ]���7����V�Ly�k^E���)xA)z�$7T���"d��r�H�רme�M~��ea}�_�5��px~P���'�5�����(�-�^�$�k@���'l�z�K�.A���JD����q�N�Qs��(�^7z���*�7���Dj�ȓ�NK�E�f�&��~UB�!�m@! �Ӓ$j��֗A�0c���D��dVj�^󦿯X��e3Y�+�B-��ϳTK@��9p|��QOZۅ���*��p�����Q i9K����&��!���w!��Q���s����,vGSB���@��7�Gxe�wA�$�nT�H��4����]��/�Պ�2%�@��Vo�����.�0�Vq���������(@g�h�r6[���ﾨ.�PD����w1�,80.����V	C,�|Vz���Y�'#h$���R��C��J�7Ԗ��
$U�d;����*�R:�	v�xi����B���Y�J��یC	H�ޙ��3�)�Hl�+@\(�����4ސv[g�䵒�5Ó���.�iMș��.Q:��Z�l33�_��Ȃ�kx�r4���4/1V�ka������+G�Yl)C�8U�:�J�Q���J�D��o�|a��R4�8��b�|&���7A-��&��pc	�p7���'�����_��0'"�v�s~��1��7d&�v��</Y���C!kF
#-����ua�/'l����X� �T�X[!twa�vkl�z]"�<tg��RZ�e�:���joH"�<.��	SN��$���N��/�Ͼ�`ژZ��#��\E�8��Y	��مfM1G!
���`����2wJ�'�&>� ֱ��y�*�j=���F�����Wᒧ/���ޑ���$|y%�z�[�Aq��w<Ua���i��wݺr-$�ɕ'�(�t�!m*'�4��!9ƾ{�&�HP�ɔMB�/kw<m-J��Iӽ�Rl�_� mF+����[P@��=�J�T���MYm+!���4��c.z�Y��o�Ks²Gw��!�! ��T�vd�_B�R̓����T�s��i-L��8��N�:�Ϩs^�� �:hy���0؞��O\n�oZ*7� ��u*ȥӊ�_�s&s��\��Km�����`ӳ?w!h����m�e7g�����L��Ov?øWBUQ)d:'	�W��T�YBj�f� �H�qo੹z���t�^T1J>�=�jWs0<�5Ŏ�Wx��-Է+�Ȯ�kP��z6^VM�?>��sV̳�D��6��3v̒?�P ���ƚ����%%��	�bK}�����%��@��ykN��	J��YS9���X���M����f������rB��P\*ݤx�SQ~?2U��t��&V�\���F���W���-�G�V )��=B�����$ǚH��Y՛�շ�k�}:P7is� 7�+"��}�
k�6+���ـXU�b��{��kE+�����\p��7&�l�^|��`��}�@Lae�\�۟7�rt���L��<����H�AEpVCh��E���D����Z�᱑PTM�m�AL��qU���&��Jt�I�gy7����H����#�]�P���x;s�ŷ�h`��^�j�.hd�����SҶy�V]�yӢt�7V P}.Er�}'�Z��l��M<r+��nʤ�� ��� I�m`����l�gm1E��d��"��\y�:��� ��f��ۘ�
cO$@k�D`����3[]D��	7#b����B��9k��w�+JbVe<���E�O��ᙈ��,��ˣ�K��Ԟn�\)D��^ϛ�a��SgF�z�D`������aְ������̊��`���
���k|'1�j+��&�vq���4�uZ6��4�Ä�G���B��:Z��]
�zh2'�<\��O
�|z���B�"Ӑ�<k����Ձ���b��	��������+�d��?!�C	!�sb]+��s�?x�2�Yi��}X���%�)<�F�{���>g���
 }�&��g�Η��٩7���M~���Ok�yE'm�'��G{	bB�1 �H'c��j �5h����c}+�MѾ�R�ׂ���y�D;���l1bKH���+]���S�!Cكx�g΄E�auGqT�W>�ɽ<E� �U����X�S+e܄�n=��9���0F.�ޟp?����G>��E9�����"���O����2�ȈCp���p�E�)	�	�����r�b�_؉5��������A�K�$B,� U�+M���{bk9~�_�2��-�/׽�]`��1�'�,���n������ey`ㅿ��5lSf�/
�;�,A��#+�Š���S��Ҵ�o����ޠ��V�P���5��&�������*�_�[�E��Q�[����8�5�)��4�Q��V�'[�02w#���#i�= ���T/�zk��q]ޝ�RD,j1A�HEH_ټdt	b�/��	�&2~p�\%���s�;�َ�����@�T7HT鷴xc1�����t؊�~A��kF��.�8�d$��G�b\�B	�a�m|�	g���n�`j��?�+�d�:Mϐ<����#
��tQ����iɜ�(11��7�j׫5�>T�{V<������t[o<]���뺍���	a���%fM��m ߳\�Lflo��OLV��!�@ab4��N��m�)u-5��O�"!q��{�f��=�*/���na��+>��\ L]Z�ȩ��Q������I����o0�Z:�{Zh������ɾ;z�Q���o�uw�7Q�`��:|�C��}�ހ<�f/Q��.����` m�	�/�4YӺ�/�@��{
vI��jRʭ��ˠ���/�+�J^᰸^�^ߨ�Si�4eG��	�
Ao,��ð~���-��`	99ExeWrh�T��|h0���d/���ᆃG�"E�9̓��8n^����&JH���)ޏ^��sḋ�YF��׀ޠ�5�O��
�m�y��gv%�S�CG#�v�&�V(�
)�{��o<� E�P���|2���
}��^:;c�V�����Q�6��A�ЯSG�汴M]v!�L�6�BC����^BD v��N�0�^��1��-��q���N{��W�B���u��WV�t񠩵�M�ST5�5�7�{�K�{�Z^���[&?@�u���s�� "��J`�XV]���FE�'��jdL��u�|����JE6/�Sy(�ѐg�R�ʆ�rY���Z� �^h�m∱���R'�]2��KC�Q��x��H���u��o�Z$��zN� +�Z�U���5�3�!l5�����z��j7�w~��&�5���c5E~��#Ҭ�a�-H}QK ��+C�-�p�)���s0����p͜�"
Q.`~t�Q�6,�mC!�����{���L<�G���������Na�� 9�#"{��0LQ&v�5k���#w�𼟤=1e,�=.�Ď6Ͳ��p�p����W�������㇮��w��9Bp���WI7pP��ώ���K� ��H.�`X���2��+C0-4
��Dn�)��Ѿ�Y�¡G�4���5F��S��P~���dZ������*8�������R�T�;���Ui�̠m
c��Q�0^!���xDF[�6������2dJ@�5�6��Cq�����3��ԅ��k��������W�U}�iز��л�r#�����b0��PӺʄ��7݌F��-9'�u�r��7��E<%�D���,e���/:[�:W��e�S�8�k9�Ђ��@_3��s8C:�ʭ��?��8l�B@|8�@��h���@yQ�Ǭ�H�&c�����U�l�2_A�[lkp��H(]_>��\'V��ozt�CZ�������mtk��Bh���6�dOw���'K_�����[��=#�`�P\c����d4Ȳ%��Vԡ ���~�`�����i�;g9�b@Tl�c�lv[w�s`Nz�ґV�v�;҆�N�"K�G������-� ��k���r�&f�{w6����8��W2��V9�"�y�P�ݻ�a|˟�FV��Q,Mx���a��G��yx�k���ޤ��,��jJ�J�x��B!�ㅊ�v����ۭ~|)�U:�}�<�ǳ��Qo����d�7���R�u�; �;y��"�x$0�>��Կg���������
`�^0|���;Q��$�:�0��*(X^�X��f��9}�3�����[���j%}݃����L]����F���bh��"u�g��m��!M=�4����7%�V�����^�t̜w�8�wJϗ�y��{+]�}WQ�T�T�T��Tu�(+_Ve≨pπ�Y?�cv�GG�V��y2�ym�d�����x�өZ:� ���qޑ�vB�j$R'sϽJ䷽����lR\����>g ��5/�2G^M����i)F��a��2���+K�&$ɘY��;�������(�b�L��E�G�"�g"5�C�%���׈u'H��γo�"��`9j�ı����|}�RX ��[�z�]60>p2켦�I�d ��g�m��iy_1�R���<����VcUElsws����/�1����7�Aͥpo����a geq���o �]�E�/DHDmj�堿����'ݻ��$�w#>�� <oS	W�7��X�|�v�{��v�����f��-s��׿9�[	��(&'x��01MO���>R�{�n�##F��s��d�ԕ��Rq�E�}�cN���;4�44����#���'�y-E��#|�����<�p�3��6�% 
��OL-(~ Ì�7���B�<��E����:�ʊi�����z!�� ����6��6���|���r�m��rO�l���h��AN`��<��Lj.�Ԑ[�r�nÉ���I*�ct��9�j����9��  �(����٭�dk���\*���������형�{���_L兀v��˩,��A��G���oO��XVoi�P���+�H���]���������Mm-@�/r���$.�q���M��T�d� �#e�*�&��]զ�2q13&���=<�h���Fq���9R��w�áfm�/�$�Ph�ra��h}����)�´���mK����ޛg����3�
B>������E��A��b5���e�|�uR�ً�j!�6���bN;1��U�W��[�;��7t�S�E��u儨hj�7<?���m#�T<�ȭW�$��p6�N��P��F�*|��Oܭ���'�������4<��jU#��A���gE�j)���ث�Z����уp/�78ܶK�h�(���ԗ���Xs���NY�`zO1��g�2L���� X�V�5oI�����k�4���ׂ�o_G&>�������K�^{�~�ۓ�}���=
�����n�Eh��~nR�,��|՜���Nn�g'�X{o_C�����U|tj�sώ�|j�Fәzto�*�O_�t���Y��m���Գ�4��I�X�D
GnB�?�oyp���u���w�.H����)��I�gYdC@��f0T^s��M�� �5cvD&�1�U-o����yyC��x���d��nTJ�)�i)H�+WV<�_8$�϶�Zc��;l\Z�(��Ql�0�e>��x�\V��#�����6�1 +�6;*��#����ͩ���$��@=���zz9cD�!Y��0����%��
0���6�Z�&��-r�o.s�ŷ
�C^[ՃZ�a��Wg����4,��ac_n������'�L�MW�����g;S��găec6��R>���ߦ],=��卷T�=T<��f0�j�k���������ܾ
��/pٛ�'z�PE2v�����[�Q�p�8&?�H�m�T�����m�d�c5S{+���*_˩��^�h��r�)��[���� iw03f�x7����Ma�An}��'�u�s���%��f��7+3��hL�/�g��%퐡�����;n�{?4����K�2��~M߷��ʇ��sؗ-%�0�tN�9��d`/x��.HX�1z��W~���e���k�<u)�Ca:B|~�?R	*�#��ί�^}=׶[�+��ٍ� ��+LɅ����V��A\e-f��Ȅ�G9j�%���m Arr3$�e�ܳ�8�L#)�c�Ɲ?����$��O�wiR�Rk��,]2b��+��b���O����yFOX)z�󛏶��+n��=��(0�׃��[E���i�K"~X�����t& �.�����M�Iګ��0��� 9��2cS��N�.���.S��RQ-+�P!�ı7�5.�~e�~�%��ojVt��9�n��R��{o6�+��^C����-)(���V�9�(Q�l���zcj�W
dEߜ'�@D��Z����9Di�'������%/tH�--Zky�x���z�z����Zl�lq��.nXX�%��]��r/��a�U���ԧ'��Z�&����5��������S+|�����%$�6ୄ.Y���#
@�A491���=g��)����C�ez���wW�! ���z+�(�U�@���X�sáYP5 ���M(q�I�!�h�I6�-���V@�t�+`��d��r\��k�l�
�ӄ�,B}��)ԠB(�o4O̖� s�v�-QKz���Λ`x�E��T�4*O��A�'��Z��`ib'u��jr�*Z
ip�Tr�׾�P�GO��,_�G┣?�2޼"Պ�u�6qw�g��~��?j�j&�66�Z�p�b�{E�Q=̥�������S��{�ٴ�x�u������0{h[�B�$�bV	{�YLm�p�������-�M3Bw��r�@��d:��6Or	��O���R�8A���)�W_���]����)�]����� v�C�<y����Ў��4�o���rn����=>M��9��/��L?���蒟�!]m��f�K�����<��Ћk�P�=ݖ�rMA!o�幗�!V��H7��~�F��A3����A~nV�J�9������(u�0�P������t�2���`/�L�C .J�-U�6�D6s&[4��T�����'ݳ}�i�Ԩ�o8�Uz�2
X�#Q<����y&$|/��&Ï�ƃ\s�e2�A�l��ܐ��J�����d����3��r��a��-8�Xd��C�S�^-���g�o�]��U.�k��A��ّ�KЯ��'���ev�J SֵL��Z��mO2�Q^O�h��8!���8Զ6�B����6��mg0��]��PRa?�K�O�vwl���,����}s/!Z
�O���I��_�_�/�H�b��*ng���F���8h��q5��l�-4��4��Q�jVNYbQ0���E)����y�S�V}��@�1�c^�*���0����[�`��㺞^α��w�c�a!GWᓍڗt^�����¢�Ѩ8���#��yD���>���CWߗZ����ԭbJ���'afV�ʙfM��u@�c�~ Y,�`���v7I��t�|�>3���j0_Tӻ<@܆�6}��Qh��q�������B?˝y�������-Hl���9{��2��;�'@9����������j>����^u����M�^6#��{�U[L���>:AV�fR�˗!�3Z�x���/0�<��:5F�Z��Y�6�̠�zA'�K���'2��>�k.ݓፅV8xeլ��p*�p���~�O6S�+C�/~{+�a۴�S^��%�|�C�����-�Zv�:k)�go�'��N^
����::�#D)F�J���g�����q ����]�3 D��~��iLK��Ñ�j��6�!����:M��(�G�9�7�U����	v��Cē��L�޲��yo�w�����Kُ
���{2�_�����X�]0@��	+X��M����wOԺ* �q�m��qW���-��Q,G>�����XĄ<2R��B�%�x��Q*��������;M��|���u�=bL	V^��]E) A���X�js�1��d�P�mB�\�������J� r��Ҝ���4�g�e�f���./چ��ҭ�`u�ɳЀ��C'��Sl.����O	0��n(�@D���BJD����\��#%�%ҍ��t�!���x
�DG�Z�P�{h`�>){�_����qR�Y��v��3tpf���p���9�l�%N�m��=I�dA��]F/��Jo�����ʱsHn�o�ʰt�J��\T�բ��8j��
Ь���U9ޓTތ�+S�<���;�H�*!���V�>\O_��<s�ygmXck�}�� *��� ����}Ӿ��(�`�KԔ� [@��ؔXn��W��k`��f�kRM�K:���������t3�QD�i�u�!��lE0����zt<e� A	�6.-'l_9m�q&�/F#���?�R��^EUg�7��7Q=��kζ,�q�QE��q����� �^KQ?t�7��Ÿ7����JD��Y�i(G��}r�h�E�B�Fఏ�a�7�/]��b�,�3×$B	�C�07D�|þQ@�L$�.�sgHc`����
t�"�)�:P��b��*P�B0u�%������ 0��/xU]C�=m"�1�5q�w��{6��RY��Ck�����TS\��Ǳ�+��R�������}>�w ZW y���1/FR	)þ#����}��[
H�Q��ksf�&d��j3���`���W��SO�'s&���Ϯ��Z�n����j�uh4�>��j�hV���Ѽw/�ę�d�f��Q�R6h�m�h[�S�<z
c�=0��k��4g�c|H'�j�>���V��.Gy�h�w�!�	#:!��/��d;}�LE����n���R��ٝ-��.��q4�l�����^���ڤ,�8Q LJ�mqu���P�a��r6��ዽ���~ųjp�SfD��azH,iQ���n��c��IK�4��f�]P�T��o�Dq���-���ʸ%���c]�{z����Ml���X�B"n�ta+x��a�lݷ�oU��f t�dEB��]�����2�u&Z�E�Pr�����H-f� �4�^Ɂ��;%h�Z7;D�LzhxYov�,1�݆���~7����Do�n
8C���l�W�}&>=O���g+Vr�h�ݪ���4�J(SoLG�#i:o5�3/����k3
�����Ґ38m��=o�h�݈�<l>[�2�;���%D'a��H��F4N/N��� ��$��n����ؗ�����^���xN�e�]�[J�\�˷�{��W[�m7�����0�o.���TlD
p���^�ym:Ԇ�ۄs:�i�\�X���HN�	$k5Γ8�"��!C�[�q�c��V0 PY�'�r�K��KTL�#^1�/�!\3e�	�+G��E� ��Y���6�{�R�d��yo�@�&�L��>U�ך�gA�+�Y�{ 9ҵک��w�s���6Y��u"�Z�XB¹��]�)u��< 嚺�X���wd���>|�K^\2#T������p��/�SDZ~g�`��5=uٹEH	�,dvTg�C���S�(�q��M�~���xѤQ�~���	1��aM����������S[&�L�F��2s~
x�yPs���u-�;	��xh��s�7Y&]�q��z>s��'�:����7�#ݿ(��|`��V(�����%+<@��.��Nb�~��O��&��y�7�zV�m�c��Pf,\�a/�ލAN �w_f��и89����s��)�岔&�U��kQ`$�y����w������AJS���J|��?�^CiVQ���0���_@�H��ܢ6I��{x���Q*t��
,G�=���<��%�Z�UK�sKXԏ s�vMM��zL��I��=A(�X'3W��2�-�l�/�K��>BA�IVq�]%&Ye�F6c��7�tR���D��h��E~�p�o*��4��%)o���)N{�k$(f*"_�?��z�1eV���������{���:w����y.Q�����9��L[~[Q�^��!�R�m8?�n�b+\���s�IPJ4�?�B����n����R��c�Gc��ri�?,���E�{� ߫XW8]��ַxq�.�7��&@�>K�/�E��f�}S7�ɿO�\�>k�s"��`��UX����y���"aR�����кK����/�/�wd��CDM�����a�[K�\���������}��g�0Em�S5�*�5ș��86y�9\��@� @�d49$�o�r�Qeu<	J/��y�:�V��!�F���"d�0AkO�cQ���3�Ѥ�:�^q�aUH��X���4CM͊1��$Ԉ�_w1�_�r܅�Nb��ޗ9?�W�c'�Ǥ�M�����3.!��z��.�M� �X��K]��w ;` ���K�._�2 �ӥ���9103rP����������nV����@����M�P��%�!�d��`.֣�W�-��ͫ��ï������]tM�LL(���u�!������[�KUD�1)��\!�e�y{��X�<e}om`�V� �4,��,�%d�J�����<�8�=�Ǿ�.Z2a��I��!C����ǻ0��w���[U�R���zVS&@s�ެ[�b��JI��֔����J�����;��M��̸`n��#�h�2�ʿ����O3������h�4c,�>!�y�;[�V8�YQ�&���v�ǫ�f6�����)VIK9�H�k��4�E��!��ǹ[�f(4}����?��0���G���$rI�0p���I)Xz� a��:R�jR�ˈ�;��ݨa�7[�����N�RHV�΍�� ��6��;B�9��|�鞐_uto�B`s����K:
�Q(#��V)C���<,++3Ģ���'�B�*8l�<�����p��*�Τ�Ks�;�������v0�5�{
�ОL7����y�D�]�����"�o�7�_wDk:V�!,,/$�P��<���s�ļ� 3�$U�AYiƖb��ͼ��S�0���Ma��~\��f\�9R��V��(Z������dL�Ĺ2�0�|��,y˴�����M՛�b	���Q�-ظ��vSg��2zd�\��=wi ��ى�U�F��Aģ� �o�/^�Y^sv0���
�s�ըk��dMr�]�8����<{��"�7�+�_'��7T����]�Qs����!�S���Y�!*w&��b�KƔ�뚺j�N�4�K�I����i�2X��J�9T�nЃ��k�%�5�Ɣ�v1�8�����B(&hN^7�q���7���7=�l$E��-V�~t�$nP�낗^������?hFR�j=���~�� ۔T��K����0#��&g�0`_ɖ�I�SЧ�Q;��N�w�ڶ y���Q����t�}��]���S��J��/�<3�*�@!�Q�r���9�bSw}.�£v�u�g�����^�icz xd=6��D�z��0�V�i�(�[�Przu�����D'陫@vAFێg,��E�ّ�Ej�@�*ǡ
:��`=�H<�S۪�5�?z�� G�y�.-�� �@��lw2y�?��YY�f�7`/3h�n6qY} ����U���:lԯwh�Sd��JI����@�����s�)NE�-2�������.W.��5_S�4�Бzkb!Iο]��i}���⊜��r9�0뗑
Y�7I�2Z�4gO�/�瑭�9�\�� �Am��+Dv����q�{���8/���u#A�6�Цy���z,/É�ε����ʹ,o���B�wY����, ����G΂�Q�Tk �#�5[x�3|�,u���p�E�m��tόs��~	4�^�����<���e�ǲ����`��F<m`p[�ai8�2��InO�Rv!cIs�p�D��H̊��loxo�}��9�F.~����8�gM}�'(�ϥ�4}�����YI���k{yc�8�;�K�E�S�:$�X;l����`l���R�
	�hZ�^��"�	�QH������5g:��5��y�M,ۇ`䗍hM�k	AX8����:>%T`���.�M-�E�Hkn��;WoP�����K��,�%��m_��f .�w҃��S�g��e�if�v���uh�C��!�f�V�i�ꬅE+�&�d-�PS�03�[`�Z-P���^�>�{Ab.��C��	���{�B�p���m���w��O��~���7��0��(v�$������"r�����Q�Y:���@�'�~dc;I���:I*�U�K�~0�$�%�F"R4D�dA��|8ߑ����<�O��SBC�4�.��:�
�:��#
��cvs'[���n1��m���&�CRgX)��d>�I�{�8u�#�/��D�F��+�,�]��V�2Q���l$O�p� $W�D�@�]�6�����TI�U?Fȥ�/(��ޚ���z�:��ރnC�M��^^�ow�I~%uuX\*7K\fʫ�o�9X)H	��y�)�a#.��i�!�+3+��K ¨��6��
���J���������Hw��2��s��̣9���P3�gwmY��T�ߣ9�s���#���NM���XA���5'2_�ՠ�A��ԃ/��{�H$�u�Fx��Z������s��ݝ��`��:�7d+*����DUs�n�}E�c	f%h��
�	�G��6�xG��C���e*RmS\k�o�+Y�[���+�q�c��t�}6�'fi��ύ�\�Tx��ȴ�X���1)3^�ϛ�7E���LF�F걍���F�D�>ݖ2�@岩��ۇ"����C�����}D�=����~���_��j��0�g�,�Xz:E����,9Nuh�7��7�c�j�T{�DA��Y.�,�/�Ī"{�@��M��J�ދ��;z��C���m�w�8$��y	�@�uYH�k��b�W���<
�ƶ��qL�^��u�y�~�Z6Y3E�d#H��쇧hJ}�}4��flA8g.8�����mը���Ut�hB��g��腭���QCU�݂��ޤ��Urd�}�Z'_���]q�p�_gn��~�E˝��%NR)�����*������w�����
�Щ�P뵯_G7�ܢ��F���No_�%��(���c��@&�yL�a2ZH����!�����G��E�+�ð�۰d������+�N�?�c�*��^ ��x�����[�[�u"߉����,9u�4vN���
͐&�*!3�vH(�y��W��k�9FZOտ�/CU��C4�K��l�� ��eh�u<��Tr�̸P�)��-Jo��̜(��ŽVwF�Oqf`���9�F�&6��d��HcXg\⤨l�ʯ���?+,k�����R�J�+Yr�XUy;ȹ3k�9�(�߇*a�~H?����+d�����jG�W���;�	j�#�4L`-ݤ�=���@���J��>x5[W��<�@�*�A����ʋ�&��d$��d�ak,�M&�e�m(N9%y*v�҉��!_(�!���p��{�zH�S��*��o"�9:ϲ=%D�D"��.Q���J���r5[b���į�أ�aF
'H5(�=@�w�c��:d՜F�TUٲ��sg0ng�d���jk� ���?�c�1���&{�!L����/�˰L��vBL&T��ќ_��N
�^�
^K�S��hrn@�T��J�_�)��Y�T����G��F��I�{"�v=x�����.���h_���ut+�HR��z�k���k][r�|��7���*�m�����⹃ǥv��U�5H������C�J�`}�Q�K�&@��EQ'�*xv�{Y�T'-��*��o��4�Rd�=��	Oas�iy����^|�I���,oz������j�5��B��W}OR���i�w�|;��q���/D�7~����S�M!��h ��M4��9�������v�=�`��b�śY�0}Q�s�tWR�hQWF犵� ?,��݆~�(��i�k���4�{�g���c�>�x3���镛�B�5:v�L#� �c}���`3���c ����Df�`0���H2B���\��1��)�_�Ɉ�K ���N�A��*{F`N��1JҘ���ϮQRI��>������>%R�S;?�������f�V�������W��;u��^��|��H�9��ٍ�����3ªU�؁3|�'`x�M��S@MN]�[���t�5�����<+�{����bLT�]�]��2b��(t<��J�wM��N��{��I�7��q���N�����-(Ϝ��0��(�"�R�G��zȂ�Vn@uDH�5̔�z�4��Aɩ��vy��_���
���p����Ţ��];��k��̭@S�� k%>�ØksE�4�$���V�e�W��;�7��NA�͈���bJڮ�k�_�(R��!���H��z#���6�����/޲i�C���%��>�4����󺶖v��I��i��%���Fm4��_:K�w$�N������w�]xB��&��{�Ym�N:E��
 ݑ�T���j�ol*u\y؞p��9�F
� �o�MB<]xM}j��.:�W�c���,o��$w�Bgne�L�
��Y ���y���o5}�2��[1'��{�<HT7f�d���[�h�XR���	��7Z���O5-k�z�����DP!��Ŋ��(�8��܋��ו�wl��ŧ/|��Ӫ$���i��L���䀇B���yEtp�0�਀��Yn&�f]��dd�-�t�!�;9�0���?�p����V��d��;T�����iӞ?���9c]�VQ�Ym�D{umj��O[����#�ԕC�����E��߄Ȑ��*��f��6�k�-��سK]���˕�Hҥ�Mx=�n�Z�0�IMo��* �"NxL�,�C�s.��rp p(\�T⇔�N�S�<eA߸;c,���҃���*��Y,�F���riT�"�_�;TOh\��d
;�QS�J81M���ľ��xu��Ȥ8:e�
��F��N���qaa��xz��Q���k!d��u��K��M��`U�@�7��>�����MO�=�L�6�"�T�I5ՠy��G��Gx{��7�X\����fE>ԙt�]�͈	'��};f��*�n��¬�l��eN��N5ְ2_3��
�����`�]#?�[U�be���p�_�������x���d�jH�^�񘭠��{O��&��j�,�Y^|�zb�{X�k��~i��q$	U3;_���)��w�/���|6fc��w���K�iz�ic�&!�J�X�{��%C�C��H�!.���ݠ������a��>r���]#�Fr�	9ۉ�#g3�x%����Q��9��/��MO��.E`��#,�w4��L��j��0Iw�Q٫C�j����p�Y�SLo����d���N�޹b�ɭ�[�3�z��36�z�*�}�J�D]7�3g��&*}�)�+��G����DG>�6c�O�#5\��H˚��/�ܜ��6�l�P]���䔓���{J�uId�������G�Tb�˷��\��:�������(
�&���F���?�t0#[_�q���"g<�h���%�*�m�	�C���u*ݎ�dm��~�i�9-��/�F���2D���ک�8��:3A���zs�_��ѻ����ͼ|kt~7��p��"#��^Z�����lk�,Q{�{WR�Tc����>&����L�Vg%gE�Wd��7�4��%)�V�~�k�n���]ޟd�&�z���v��֟�M!�&��,8�`K����W��Ёy�*�T���h�;x���~�N�����kݾ��LV� ���'?	�a��������ʉP����ٷFR\�7��"Rx�����7��������_JK�# ��(S��V����^�'e筕Hr{��Ͻ�k�FT���9L�n�hƫ�o2�)�0Fu|tq��9�Q΁���@���u��*%�.ͮ�C�?&]�	ou�*\�_ws�'g���ߛW�p�ՕH���>�^vZ1�_[wԊIZ/��� �/�����I�Zv�����%y��h ?xd���MH�݋.+��IG!07rE �v���� �ܲ�z^K����W>j����b�ZF�����L�ġ0�O/�/#S�Ղ�Qg�+���d�P��K��GkV=�)������_|�y��3V��d�o�nY��fH����
Ʉ_ �s�f�.-�_�Qz�SzX��7�|�q�+�&��u�⦆_3��y���R�_>��G����N�Q��-�6�>�����N>�����,��(gH*?�C��'��a��l	Q&��>uE`�%�s�Z����ɵ�-�r��@��ˢ�P�}���aߺ��6!�V�Q���@�Q?b𬦋�lF��
ڑ*��ܼ�@����\���:�w;G���2�ѿ"��k��4��>Q��tqV���������k�b��=�I�����E�H�l�6֋G���\=����F�����&�
Ȅ.��w�"e����p������������2Z-�+�w�9K�g�����	O���/� r�=�=�z҆џ�0���lAzo
S����٥����:�`(��
+���R����*����F����k$������j�v��K�}��2r`�!+�w���<Y``�t���l�D$)�F;@#c֤����Y�p�	���%U�L����C�!=҂3�Y���d-��J�:}�d�NY��ʞn���x��5��K�i�G�:@�qߑ<�����4���)��i�i�5�D&@7t�Dv��i���sZ���V?�3���X����@�~�-�a�X�&}���5�4���C�հSTj%�c�gDl-l���"2�0Y��*�]�暴e�&lӑ��̔�.�ӣ�C|{���x���g�`@��!ׂ��6ϝp�>���NO�N�@gJ��<�:�!���o<�򇹨��)I<�d��#����KeQg�K����T���$��F~c#�ײ�z*���s�U5]�$ޗ�:3�o:�';���&!BDMZ)lg�������ow����ʯ����#%�����9<�L�'��1Eo~Ȕ��3@ʰ��7;�+w��]�ݟ�����T�PEM��g�BP
�ޅ�kk�`q�����E
.oK_�2�a�8E�� }�m5aG4H3��v�:F�ԗ��ʴ+)��ր���Q��B\���܂AGg��*�~��3��1�; ��gP5҃9ߚp,J�㒈]���>ԍ<M�Ҥ��L$�����ǖv����ɇݭ�Ќ�����A�j1mIߵ7F�3���4Dޙ�Ձ�$W�nvO�sH*$��7���؈�p�'����&@q�z�$8$(�9� }a�ǄO���L�Ὸ/��p%*%y�q�H6<�s��{ʩ��J�^��Ve���o��bf,]S\�o4��7����rʺ������73k^�uYxޯҤi��ϋSߠm�<��v�M��b�5���ۤ��˗�������*��|� yHs�U��04Ҥ����o*���C71��aN╖����WfNd�Ŗ�g�I�c\
�7���Āq�f�;ЊY�u��r��p�� 7��Ξ�� �ʔ��m��:%5�+��97Դ~�q�ϲ8���W���ۖ��ڤmo��"�|RE��O��6��ߘ+}�a/(q��c_�
}[]�&�gR�����T(&;'$&o�j�n��`=�6����M��2�BK�vi�yiK�����CRj��5�#fD�h�,K�	_�` �P��&x$/�~~5%�	ˇ�ؓZ�]�]�&Ie���l/(������J�h"�c3��ٌ14�� �{��1��J��Sg�$�D&�Q'�gaJ�5N�ON9����BR�X&6�F���J�:�,�u�{�]=\T2��R]xCXu�����NU;sMv�,HN\˭��B;:^��&�̨�	���.Y�L\�w��A����o7��:tz?:D)K�	1���I$[��V"��[ZnY�"G&�*O�R�8Ӊi��Fq�q�uK�C��U��SA��0�v"��H����r)5���`���Dg$_f�ȑcK��$�	��(�xx�M�F�ߔ�"T��T���"e��|#'/��R�]_3M�Q��3�!1�~���=�!��X����(/u�����6����>�kN��=N�u/W\6�C=p���l�Uk�&Vς�H�dʚN2UV�q��P��T)7e��0�m�
�+��Ӑ#��c�懬2^Oy����0�i�R�C�����k��*ӻ}os�IE���&p0$V/Kk`�����%�#��QJ̶X|�0�B(�a�[ٶ��ſ�����ꮜeN�;�'��w21]��e��S4��mH~P��d
����,��2S`�X�)��q>b8ߙ�g2P��O��4{��O�EN�G�6�`ڍ}��G�䱗�2�]~M�)��`;���4���ZB����a����zg�P���襀�������,>�i�C���4�F�J��>/⽙������ނТ1�l��$&}#�&� ����v;?���~��f|��MA7glY�,F.
]Q���ЯSg��Ml�
�m�����Gb���bQ�:%�tv��N�ٍ�P7��<�k��n�ҭ	��z����,^�[dW$j�m'!> ��s���ܞ�9�ץ���L3s0�; l"��;�|+��-�(��i��M���d8�%���֘�x�p�1�G�%Vѡ�K��!~��Ea����ɵ�c|��M��Y�L���үW���^~sZ����}cV(�`sC<E��Hh7�����o�/�d(��0�2�i�
��>[ͤU�Ϝ��H���e0�$T���9ײ.j��!�q��5��ū��{������;��oi�Ae��)�m��n�����x����!�D b������o2��)�5�Y�O�M%5�µϛš�Qn�w^u���G�"b�E�Q��{�+{m<����M��]	��(������ɼ6<��F��<(�����j�`�s�r?clF�e#���+�{�$�VzW��`0�e�Ϝ?f?~�k�@���-W� @J>�@�x�,�؁�d7�a?�k���{��N�칹i�ŶJlK��[�>�a00=� yH
Ou"��Fw8)�Y�Lg,�5s�f�,zT�)*����E?����ЬM�����.K�0��xihxz	�Q��e|�Yא���w)��NZus!���ʷHʻ�H��?�^�	�W]�H��fP��e��,-PW��h�����k�7�Gb��Pq�.����]�7�Z���R;1����\���|�B�rؒ��$}A6��_�NA���#Jz�݉�^�t�m.� ��_J�Ѵ�Lߵ$�&wR�:�+u1��x)Ao�7�}AF�k� 
��������Gl�2�g��{�vMfr�X�w�y6}�ǀ��'��@�>��zҤ�e�hC۴�v����p�EO�Q5�7=Bl��6b$r_ V�2ڨy&���J�҈�U����Hi+���H�u�/��ƣ)Y2�_q�5V!���.:p�����	�.x�EA�O�!l6��q�Ճ���W.��A`�C�o��'ѓ#`a���Ot��I���
��v6�`S<��X8�"Ns=�<�M�!:��� �Ҋ����[B��jfV�(��6L2�,�J�s��ډO�6���K{?!$�}�uz���g�X����'�M�1'A@y�Ά� ��qy��KejNb��\vp�A�oL7JW�d�=�.��#qy�q<���t���O/U-o�#U�-��.�����V�1�%u��;��z�,����v��@�<��/�s��C�[��(��3�fN��Es�� ��~��|�ؓL@5����T~�7��:J�^��>s�H��u�CP��������}�L�}���%��3�I��m� ������_��b@�<-5�C��.\wM�9��W�O�B��+�*^f��%؇������s����tBxz�@s�hV�y��dI1������PY���p4�Aq;�����CX=��)h�����5�9L6O?���+&=��Y3�d��Zȁ�y��vu��i�$Ҙ9�8�������t�}MiN �����$NW 8G!�\��OqC\�w�u�if�|�ğL
7���f
���_�0������+�c`12%&{�Ps��	��ܻ�:A��� =��!s��c5��Rd� O4���#<�Lyj�vPz���L�c[���ߺ��2�(D�t��kދ�=o?��*�8䭮�I��S�{(�����F�Py��T١��C�K2�gx� �M"��F-٬O�����Ά{���)��\��Jk&q��e�*��f3�~*;�) ���O¢����J��z(�Ϟ�#�?�*��M�TS�8�d�74_��Zz�}��|l���Yd.�D�`ހ����M����~�A�g!~�ʠ+�M���l1J�M���u��P����-&s���#ݨ�KM�����s����a?� w��f�,#�P��f���n�x�(h���Q�r� ��Hj��4�Zu�m����<(�#.��Ӆ�uxCb�!��Dmzw���:t�J��P]㝷Pe��A����o��|������w&���Gdi�I������nc^#�s`���@�j�a�����=�%]NΉ�3��L?�n��Ssߙлjt���"Ж4��j]
�R�HK�$o�w�N�ii\�� �(����Bl�L�rJ��ę�0�nl�
����:v�bG@��'�86T�0���k#si�����쁹0���P�DÌ����%���W�}*Zcp\vJs���O��x��{���D-A��|�M����M�S��rs��\�T�IΌz"�M]��a��Ϡp�!j5D�-4^֘��伖�2d��Y�	3ƛ�f�a�@:y�}R�s��N{�2ڜ�
aGd���3]%�q+��}S��Z ��ਅU������ �WشGt ��.8��7��tu�<�o�����Ȑj�	ԆGGn���̔��E_���HaЇ�:����جئ1�)���^��}���	r�GR;.�Hk���)�7�cϯ[�clIO�m�1~א�ܝ� v�� c&)/kE4����:e�g�Va&n&�}���+���!o��Z}�c�rx\S ��C�� 5}'�)�$�v�㾨���u@I4�7�s����z4��݊�Q=��Ϝ���b�ː�K�THl77��q�Jb�q��8�)����эwc�5v;�JW�n�w)y��HKĸVo�+���>�&�1���w����FU��8� ��bk�G��}}�=E�R��S���϶v#ni���oUB�.n�/-As���a"� kzU��n�8W���$�ӡ��U/��5{�0�RT�<��û���- Ʌ˦e���|
v"�-�ZlA�(��./%�[�Q6���w&�i*4��70P\{��q�.�} Sme�n��s�y�0��15�9���"z���Jyaw�x��9��&�1��E�7=�����]DCjg��i��8;���t�n��C��5��갭N�C����={�0'!�)��&OO_Ů3��@2��BAd���?�)[^��\,6>\e�,�P�N�c4�J	��Ib�Gc��7�B�G�N5�X��5��*�J��͓����+�q��!y����B�z���� �����W땍Hʁ�����%@
jm$U�Y�ꬶ�YI_�S
w���ļ�!,����x�v�˘�"���R���j���d��m�zU���j�0{���Z�ixf��[�?됛�k�ƨ�<�'�k����U�}�N|�����[�S�3W)��Q���n����-]���u}��=>y�¢y�cet:O�B��N�����?�`^p̒y����Gw���o��={G�/TV�Kh�%N�`�f����P����}D7u+y/4�p��d�W�+����؄��K��ȤRglㆇd���g"���镪��H}��t�N�� ��E���(J��p�x��M9%Q#�H�¨Z��
 ��_��̓�X����&���(��h��95̙y�X'�r�3���)���s22�O�JC5�c|�x��H��.6���td!
 ��?��$�����^���-���U��;�s/���R����i�-/���5=Ɵ��/L��	�,=��n�Ѹ4xdsvt�Vfk�	�j�Gw�%��}T��Q�H��s(54��Ou �.}�7�$��P��ԉ�9��j�����W���ɔ��!jJa���It
a���U���)RV|{��E%a=�z]��:�����A}g:,�?<�\�0-��xO�n�
%Qʫ`'�8K�'�r7�L3���p_�<�.����/k�z�øϏA��m�o	�k�������Q:�3>��j�yjl�t<���n[\ �Tv�����Px왑�����@�����F�W�zL��o���~�]����?;�x<_���S&x�FmL����Ӣg5�+X����������P]��~��9l9�_�i�t�^�_|�}�������gl�����D�C;�	l����tY2�ll�_�X�
m�(���9*;[���w�eC�Z'�� ?�-L�����'��������I�O���V��IL�O�R	ⷫ�B,f���R<`��Aob
����Ek�v�*U�
txԐi1-�-|<!�~Lw�1��i{6S����Hc�@=w��@�B���.H�yHTX��D}�'�Ac������j#߶���]s��Ѧh%eGH|���P *���=y��W�0p�@p����kĚ���i����oրe�/�(�	� ��VRJ�l����*2��Q�I�"4Ϯ��y�x�P�e�D?}�T�p���X�v�~AA��ɾul���`S�N�iZ�ݛ���١'E��3�Cm(}��
�:�T\GT�~��m��$��ډ{�Zx�AR�J$5��GMViI�������Y�4Cy��;^�|�q��e�(��'׶��ro��|+��wOg͗d��}�ґi���9V+$����<%�w�n��ݛv;]������}�Ŷ6z&A�c���03��[�Ϧ�G�W�%�<�
Ø�����2�d��ǅ��)����`R���(���ȝ��X5�Mo	�`��d����Te8�����]��QWM��t�m�߱��YGpF{Z�ᐙ��	�Ors*�wb����=�����ɖ�5v�T��Q�U���'�"�cut��d���<��$�Z`�Y�S��\m*,��d���r�[K�0+y#]�
/��Z	��ӽ�l�΀��q����2O�6��K�^����A���#�&��XqC�����'�Z�_��k<J�%T�cN���dZ��2|�I�' �x��fێ?j��v���g�O�������Ri�2�vW&-��-c��W 4<�MAs�����~	�8ܳao`��>X�+�ۙк�jR�h츜��M%F,���P#S����`��%��k�.�)Q�����m�H -B�tn�<��|�;J �Nԁ�?Bځ� �0�߁���Ă���9)�w��r���WW�m:�r�O7����� �N-!<C�c]Ŕ6Wki�(�ol�m�Ԫظ+��$Ir�c������ś�2�I��{���~�ԩ�|�8��������"�YQ2�'͍�R��l�_4�R>�]I)8�̘�*���L������ټ�gꇑ��Kf��V��]D�t�q�I�4ҟ�/��(~�����DV���_��"(ӺҦ
����7�>����ҝ��
����LѤ�\�Ϯ f͵�Ki������r61PJ��*��:��֐j�6;��GI���3i{[`N�b]d�1�n�j0j�΄j�W)�z?S�e+�7��Q�����9�U�!�	�$
�#�H*�D-���:u�ԑKOx�pmA�3)6Rԉ%��n&6�GW9Q�4�*l�H9=qE���!���S՝���ۋq��~�����Y�h�pZJX���C	<1"��������b+��L��m;�>�(��p��^r�x���j� x�*��O��]}�;��`�'��	M�)��O.KP3�fmzv�,��ᥕ%y&Y5�d+���29���rO'��8~�/��W,����?�-����9��mO�!�b�����5��0��/* iꦡ�|��s~������$����<�&٧ۃc,��ޘA�4�/�]vie��F0q�
EN.x�3]+������n=�.%':���������)���^�8��ON_�x��t��cqB��D5�^� ��^z.�m7a ��;���| ��2�nEe��A���T:H��Ӈ0t��0�,D�`��j#�ؓC/�}q��א?���{�gUK�b��$�&�g����i,�@������ϐ|&�?��S�ː9E2��7R���n1��Y�TӄJO6rذ8KG"���d��QʿΕ�x�T@Hg�U͈�k���O4����=Oˡ�u|`���Ck�Q
��O���Kq��u.��0��D�j����}_*I�d]�Ǫw�e��ȷ���!��d<z�{�I��	X� LF&G�E��X2���@��#���3i�~Lˆ�X�x)n��k{�oIvF6�Y��S)� Ln�O,�*jwt�ZØ�}o�)���Sh�k�������iZ���{�IB��M\}*x�Z$��\��D���F�/o{���� �H�����6d�o����.[ըΜ�B��\>MLxq��a �ْm�>W�q|�:#?��K�w�P�E��,�?��Qq��ݡ�b�c&ڻ��-O�#��e�f�D�,�õ-&Af qw՝�^�o�h�t�N��ORPy4$�t���ͣ�0γ���xeP��3hh��`�,�^����i/m�)/{�W����r�#�"�v��=��d1d"*t�BtN%�_��?�������g��S]p�{�4�0� ��P)a?%���,�OeK%��N�	�7Z��������[�|�8���w�O����N���i��Či轒a|O?�򼒌���)o^\��+wBSӄ�ۧ�N�i+���;hw��������hL|A���L�}��1�
�2� ��@C(�\l3��)�:0Cw���^���e�5L�)���f\ƽx�H�R�m&�/  ��X�m�m�}f,��$*����c��~}#��g�?˰����6�}(��לi��P�7�'���`��;`�H�een0�#%L����C�!JA�z��E���|�g���A҅ܗ��ťa����}��1�ô4��ڶL7�oDCq�����(w�T��#���d�*�x�N �z�5ͭ���Ie^2��x���%sX��jal7Q^`8�������#�_�pݸ�;_Gp=�������V��c��a_'����=l��@E�
`o�� �~�K�Y��po+��L��/�e �����?�H�����X1{��{�b!��	t:B��QX�=�	!�m�l^̶ݮX�k��eA�rТ;]��|C}	-���n�}R�����P6�M�=p�i~��q���;�±B��_-}*��6Q�	.���άڧ��ShԵ`k6�`�:�^�g�Ԥ�Z�����$�`�u�ߘD���=�k�rhb�nj�\B���ܲ�~</�ƍҸ�1�E�z����j5n	W ��}C[&}�KG5�gRy4k���n����V���$gjX�V&o���M���"X��d/\���=G>~"�RJ��3S�cۣ�U6xVWf�I ��X���V/U"nuӪ�?���vI�L�(*,;3x���߆o+t���+K~G~�,�rH��o��~YZ������C�FC7��Kw/m��c����X�m"�'Ox�ѯ�����^�{]N��cs+��;�W�B�L@��t�*s��a�/v�R�Vm��'����L
�B8`M�eNoY}�`��s�f7�kvC�{�P��8ƍ��5E�����rzZ�V"���p;\d"�vB1y����"'��>Ph�������T��r�V�����r"���8��_���,���n�J�7�e4�9ЩV�ק�˜:�G�]"�m�Jxg��1K�V�2����l%�*�+i~�%:-��Ԗ=��^�������S&oi%bX�n�ɸ����}��_ل���9�L̒cY�u�S�zzpX��"����p��������t�1��?��2)��F
���	=�t��Q����-�3K����y;�PR"���� �?�sL��'&w�اs�+2ސf��O?�G`��"�8��N��p�k�1A��b��Rk�֕i�H�����d\ �����UJژ�Q��Hyw��e�&��8J 3(�7���3��.DC4Q��(�ې�6k��S8=r�Ft��.@E]�&.��o��"�9F/�S7�"�.Z�_a��uo���.+�P�V�U�!�[�/!�5�|,1;�6҈"0AF.���.��r(����.�]R:oZ�%�Xc$!��q���l��و�f˵/��}P�L�>0�9������~L��^�� ���|��e'����|(�S�#},ʛ!�p����$�՝��FA������[�AدNx���v���6!F�� _n���g7� �>
#�#����~�{0����֞�+��l��ij�mwKn^\1�4�E@x��ޱع>�{������}�c�������^kUx�U�p�Hz�K|�fu�t]w.������-��Z-/�2����
��,C�1���E�qװ �Uh�n[�!�K8�������*��,rvQ�7�=�<dd�?;ݲ��=��30+�
���L`5x
Xz��V�I�|�K2^�7���Ź�|� �<u�R�.���@�s��c��?�c��ˁ��� ��Һ%�Xcހ���71��D������4V�������{�E]����pc+�rnu�p���*T�y����	(�����끏,)S��2ʹ!����*c�Y�z�ul�2��z�����=Ff'��r��-�<l������*m����\���Sr'��z�0�R?	Ք*`�[K�#$��][�?���Wv���"�ذL��$�?Aש/��߁c�S���K�!䇛j�Y������v�������rd�|�)Z�f{��R��%D�C�#%����qP���1S�2�{Ѭ��_Ь��', tc�e��	V=RɆ*���i�qG�~5���rȨ�RZo��M���e�	hq�6�ó�,��쐸���� ��$�Ft����}��I	i*M�R�??�5��S,���GD��뷩�/�<��)��?Y+yM'����}N���#�+�5�� �)
�ʍ��M��&J90��M˃<W���nw�؟���Y�8�Lq���œg-���s�V8
��>+�����G��@t��V�ⲗ�J��K��Qk��T�\P���-ʴ�V~ڡt�ƃ��綴��;��x���ʎQD��6���`c뭻�B��k���HchQv�8&���+�x=�Y�x��>���%�A����T�h�<qp�3�0�9��1���I��3�i�a���9ʌ�nƇ�p����jǎ@*<�� �C���wR������Ӡ�iLR�
��Sn/k*�ː)���'{��1�|΍�����^	��v�Mr�,�
��y!�� \�pa�ëG�'�����鬰nD�d|�jK����AM���X�_�ـr}+���-�������yټ8������5e�����ߟ�ۧ�m��mz�C��ܨ�Q���������D5�á%���$^X�o6��P��rC�F��}������{ӈ�w*V�vDD.�нY�z����q��������D�g"<iꚒ-bTB��Aٰ�zC�0��@�4�SnGl�&����-Z�{M���nFa���p���D稧I��a�<�OH%+]a�$���Y��s�o�A�zR+>�Pa�|���(GFMVճ)A�?�r�2�q� ݙo?#�c��̪]�!/�?� ]Q�D[�F���j��T.N�C����B��A�|��<i@�ɞц�G���ےQ���o��:i uȃ9�o�J�ۚB�|�	(�X�=9��]ME�8J.Z< ���Q�@roE�r�R�����J��T��ۆ��5��rs�I{GO��G�ԝ
!+9��	"Q[�:Ծ�h��2(^�u�
�B_��3TR������)��+�;}�Nќ���^y �=�����ً�c�������4�aM��1܁t����9����7�.��c<3���;�h�?&�S:�z-�!�jW�S�F}tM�<�ST���!�%�UW.�I�ї��(�;�?�{E2c��"�$�*����,Yjs��>���q�m���83�#�j-G�[�������!�ԒO=\�B�	/����p�jQ�d�]ے�TPd��-�K#���=�\�ź��p�]���[%���ePxfWp�#>i��܄���̷E� fQ�[�C���*����s٣/H�^�S�D%k�Mb�Zt�M;O|,�Y�t���Ʃ�
Ǽ�:�p���HO�#�e1���|fP`>���َ'Zڈ�7^W-�˳��h��|e�l��ZȕFRW��±Ȳ�|�PJW:�@7D%��$��������}`/���`4]�6@qq�
w�{����2���y���`������=}�A�O�1��F��9��B��j��A�t�3��K���a���\��.	����\fg��wu^�c��EsK�8�$_���:;�����O<��=UR�&|��(#J��a�¸�<�;!�����}�e��(ȧ5��f���b;z�>+?*w�>�V��]�C/�� ��ʋJ�o����I�s���������O	�/qh�f�P�؞��`�y������>M6h!Jd���o���@�c�,��g����Bk�4�gP��܍�a>��8R��.6����ܥ����e
7��x� o����p<cx����W��ނ�2X6�i )��WA��g���z�(X83��^lR_徾5��o�3���guҟ���#��8?X'�	{�U%�Vq�	y~����]���80x��d�}1���t���ƴ=�2�����c���?�ҭ�
d�<����E�au�4���B�5�os��e\�2�^L��G��'e�!kg	��V9�(�rEn��j�ג+	A��*��ݘ�����Y����X%�u'Y� ���FOa+�7.=��x�?Tr�V��U?x!���3*�h�����5��!���*U<�궷�4�m�lV����%-� l��Nn�"���g6��8��`��O;�w}��V4"f5@lsD�ǝ���4ҳ�&8޻?�5��~�Q���&�v}�N��yT�w�9t���JWj����/b(O�e���K�K��?��1�*�����c��q�0-*0�ة�E*��I�$����9�C{��B} �	�	4��ydi��~�{�1л:��G������o$��� ��4	�ǤJw�t޻����z�&�, �@����':#�4F�r��i�2�b�ְK��8l���v<w�͍���6i�g}L:i�PP5�}��ѭ�I�����pȨoon�K�n��8"�l?�D����a��_Y$�;��z1#5��kZ�V�)�����^bY�3�==�@���VpFA�m�u�9����_1 .07��B����X���	9�St�b�f��G���6�\�ܴ���m�����t�PL-
�\@�dǔ�{L���mp��o^��\>$�QcvvE:��,~�����gJI������@��#�o��8ݻ�|Ly鄤��QO��H�Q��g�5���G�1������ۑ�H*2��U&��|hDs�H��{����V��l|��٘�TI7����!��LS6�2��Ίu8]�&8�����P�E��U����m	�=�����QH�O��:3B��;��� ��z	Q��b��	�I1±Q�9Co�Dʽ�Z�h�����Q������/=l�}@�뽻m�=B�[�8�P�sD>߄z9pl\��.!�;_��ņ8�m�g�>t�Ň�&�T�@�a$z�}�&�o�Di����WFc>9Z[��k L+ @z��8�{.̌�cW���q.�0/!%Ś'su�_�DJ��e���rsF���8��Q�D����qо��WP�Hbٓ��hus��n3�c��'�ĸE�����)h|_F�𧖎Gx���u!,���}=�>�0Í���ӣG���o��g����aM+;�B	 q���^C�+ţ�[���Ou�`Mo�Vo4uT]}��8m�R��%*��)��G-���O FG��B��y`;>oYY������=���"���!	��R,�3�~5����|�c�D�"�L��b��+��`������2Ă[;��`XqIl�+t�ښ��w�̜yoyRf`g^-:��VA��s�����Zԟ�{ui���g�t�l$�&G6[�Y!?��A��Z����,3DOfy�j����uWT��(���UF����O���.{������'r/��%��{$��R�gM�iz�����[��!?s�*��ѽ"��1����b�KcG��Vbx Զ|�4�Œw~���|e�|-o	G1�٢8v5�<��,�Q��.R�s����Wz7�0�B�b$��ȍ5*8�ZUuQ��[_X~�����T�P\�-C�a�v(�#+\e��X���R�P���JU0���@